module csa_tree_add_104_26_group_173_GENERIC_REAL(in_0, in_1, in_2,
     out_0);
// synthesis_equation "assign out_0 = ( $signed(in_2) + ( $signed(in_0) * $signed(in_1) )  )  ;"
  input [8:0] in_0;
  input [1:0] in_1;
  input [15:0] in_2;
  output [15:0] out_0;
  wire [8:0] in_0;
  wire [1:0] in_1;
  wire [15:0] in_2;
  wire [15:0] out_0;
  wire n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57;
  wire n_58, n_59, n_65, n_66, n_67, n_68, n_69, n_70;
  wire n_71, n_72, n_73, n_74, n_80, n_84, n_85, n_89;
  wire n_90, n_91, n_92, n_93, n_94, n_95, n_96, n_97;
  wire n_98, n_99, n_100, n_101, n_102, n_103, n_104, n_105;
  wire n_106, n_107, n_108, n_109, n_110, n_111, n_112, n_115;
  wire n_116, n_122, n_123, n_124, n_125, n_126, n_127, n_128;
  wire n_129, n_139, n_143, n_145, n_148, n_149, n_150, n_151;
  wire n_153, n_154, n_155, n_156, n_158, n_159, n_160, n_161;
  wire n_163, n_164, n_165, n_166, n_168, n_169, n_170, n_171;
  wire n_173, n_174, n_175, n_176, n_178, n_179, n_180, n_181;
  wire n_183, n_184, n_185, n_186, n_188, n_189, n_190, n_191;
  wire n_193, n_194, n_195, n_196, n_198, n_199, n_200, n_201;
  wire n_203, n_204, n_205, n_206, n_208, n_209, n_210, n_211;
  wire n_213, n_214, n_215, n_216, n_218, n_219, n_220, n_221;
  wire n_222, n_223, n_224, n_225, n_226, n_227, n_228, n_229;
  wire n_230, n_231, n_232, n_233;
  xor g3 (n_80, in_1[1], in_1[0]);
  xor g9 (n_84, in_1[1], in_0[0]);
  and g13 (n_59, in_0[0], in_1[0]);
  xor g14 (n_89, in_1[1], in_0[1]);
  nand g15 (n_90, n_89, in_1[0]);
  nand g16 (n_91, n_84, n_85);
  nand g17 (n_58, n_90, n_91);
  xor g18 (n_92, in_1[1], in_0[2]);
  nand g19 (n_93, n_92, in_1[0]);
  nand g20 (n_94, n_89, n_85);
  nand g21 (n_57, n_93, n_94);
  xor g22 (n_95, in_1[1], in_0[3]);
  nand g23 (n_96, n_95, in_1[0]);
  nand g24 (n_97, n_92, n_85);
  nand g25 (n_124, n_96, n_97);
  xor g26 (n_98, in_1[1], in_0[4]);
  nand g27 (n_99, n_98, in_1[0]);
  nand g28 (n_100, n_95, n_85);
  nand g29 (n_125, n_99, n_100);
  xor g30 (n_101, in_1[1], in_0[5]);
  nand g31 (n_102, n_101, in_1[0]);
  nand g32 (n_103, n_98, n_85);
  nand g33 (n_126, n_102, n_103);
  xor g34 (n_104, in_1[1], in_0[6]);
  nand g35 (n_105, n_104, in_1[0]);
  nand g36 (n_106, n_101, n_85);
  nand g37 (n_127, n_105, n_106);
  xor g38 (n_107, in_1[1], in_0[7]);
  nand g39 (n_108, n_107, in_1[0]);
  nand g40 (n_109, n_104, n_85);
  nand g41 (n_128, n_108, n_109);
  xor g42 (n_110, in_1[1], in_0[8]);
  nand g43 (n_111, n_110, in_1[0]);
  nand g44 (n_112, n_107, n_85);
  nand g45 (n_129, n_111, n_112);
  nand g48 (n_115, n_110, n_85);
  nand g49 (n_116, n_111, n_115);
  xor g69 (n_74, in_2[1], n_122);
  and g70 (n_123, in_2[1], n_122);
  xor g71 (n_73, in_2[2], n_123);
  and g72 (n_56, in_2[2], n_123);
  xor g73 (n_72, in_2[3], n_124);
  and g74 (n_55, in_2[3], n_124);
  xor g75 (n_71, in_2[4], n_125);
  and g76 (n_54, in_2[4], n_125);
  xor g77 (n_70, in_2[5], n_126);
  and g78 (n_53, in_2[5], n_126);
  xor g79 (n_69, in_2[6], n_127);
  and g80 (n_52, in_2[6], n_127);
  xor g81 (n_68, in_2[7], n_128);
  and g82 (n_51, in_2[7], n_128);
  xor g83 (n_67, in_2[8], n_129);
  and g84 (n_50, in_2[8], n_129);
  nand g105 (n_143, n_59, in_2[0]);
  nor g108 (n_145, n_58, n_74);
  nand g109 (n_148, n_58, n_74);
  nor g110 (n_150, n_57, n_73);
  nand g111 (n_153, n_57, n_73);
  nor g112 (n_155, n_56, n_72);
  nand g113 (n_158, n_56, n_72);
  nor g114 (n_160, n_55, n_71);
  nand g115 (n_163, n_55, n_71);
  nor g116 (n_165, n_54, n_70);
  nand g117 (n_168, n_54, n_70);
  nor g118 (n_170, n_53, n_69);
  nand g119 (n_173, n_53, n_69);
  nor g120 (n_175, n_52, n_68);
  nand g121 (n_178, n_52, n_68);
  nor g122 (n_180, n_51, n_67);
  nand g123 (n_183, n_51, n_67);
  nor g124 (n_185, n_50, n_66);
  nand g125 (n_188, n_50, n_66);
  nand g140 (n_151, n_148, n_149);
  nand g143 (n_156, n_153, n_154);
  nand g146 (n_161, n_158, n_159);
  nand g149 (n_166, n_163, n_164);
  nand g152 (n_171, n_168, n_169);
  nand g56 (n_176, n_173, n_174);
  nand g59 (n_181, n_178, n_179);
  nand g62 (n_186, n_183, n_184);
  nand g65 (n_191, n_188, n_189);
  nand g68 (n_196, n_193, n_194);
  nand g156 (n_201, n_198, n_199);
  nand g159 (n_206, n_203, n_204);
  nand g162 (n_211, n_208, n_209);
  nand g165 (n_216, n_213, n_214);
  xnor g170 (out_0[2], n_151, n_220);
  xnor g172 (out_0[3], n_156, n_221);
  xnor g174 (out_0[4], n_161, n_222);
  xnor g176 (out_0[5], n_166, n_223);
  xnor g178 (out_0[6], n_171, n_224);
  xnor g180 (out_0[7], n_176, n_225);
  xnor g182 (out_0[8], n_181, n_226);
  xnor g184 (out_0[9], n_186, n_227);
  xnor g186 (out_0[10], n_191, n_228);
  xnor g188 (out_0[11], n_196, n_229);
  xnor g190 (out_0[12], n_201, n_230);
  xnor g192 (out_0[13], n_206, n_231);
  xnor g194 (out_0[14], n_211, n_232);
  xnor g196 (out_0[15], n_216, n_233);
  xor g197 (out_0[0], in_2[0], n_59);
  and g205 (n_195, wc, in_2[11]);
  not gc (wc, in_2[10]);
  or g206 (n_198, wc0, in_2[11]);
  not gc0 (wc0, in_2[10]);
  and g207 (n_200, wc1, in_2[12]);
  not gc1 (wc1, in_2[11]);
  or g208 (n_203, wc2, in_2[12]);
  not gc2 (wc2, in_2[11]);
  and g209 (n_205, wc3, in_2[13]);
  not gc3 (wc3, in_2[12]);
  or g210 (n_208, wc4, in_2[13]);
  not gc4 (wc4, in_2[12]);
  and g211 (n_210, wc5, in_2[14]);
  not gc5 (wc5, in_2[13]);
  or g212 (n_213, wc6, in_2[14]);
  not gc6 (wc6, in_2[13]);
  and g213 (n_85, wc7, n_80);
  not gc7 (wc7, in_1[0]);
  and g215 (n_215, in_2[14], wc8);
  not gc8 (wc8, in_2[15]);
  or g216 (n_218, in_2[14], wc9);
  not gc9 (wc9, in_2[15]);
  and g217 (n_122, in_1[1], wc10);
  not gc10 (wc10, n_59);
  or g219 (n_229, wc11, n_195);
  not gc11 (wc11, n_198);
  or g220 (n_230, wc12, n_200);
  not gc12 (wc12, n_203);
  or g221 (n_231, wc13, n_205);
  not gc13 (wc13, n_208);
  or g222 (n_232, wc14, n_210);
  not gc14 (wc14, n_213);
  or g223 (n_233, wc15, n_215);
  not gc15 (wc15, n_218);
  xor g224 (n_66, n_116, in_2[9]);
  or g225 (n_139, wc16, n_116);
  not gc16 (wc16, in_2[9]);
  or g226 (n_65, in_2[9], wc17, wc18);
  not gc18 (wc18, n_116);
  not gc17 (wc17, n_139);
  or g227 (n_149, n_143, n_145);
  or g228 (n_219, wc19, n_145);
  not gc19 (wc19, n_148);
  and g229 (n_190, in_2[10], wc20);
  not gc20 (wc20, n_65);
  or g230 (n_193, in_2[10], wc21);
  not gc21 (wc21, n_65);
  xor g231 (out_0[1], n_143, n_219);
  or g232 (n_220, wc22, n_150);
  not gc22 (wc22, n_153);
  or g233 (n_221, wc23, n_155);
  not gc23 (wc23, n_158);
  or g234 (n_222, wc24, n_160);
  not gc24 (wc24, n_163);
  or g235 (n_223, wc25, n_165);
  not gc25 (wc25, n_168);
  or g236 (n_224, wc26, n_170);
  not gc26 (wc26, n_173);
  or g237 (n_225, wc27, n_175);
  not gc27 (wc27, n_178);
  or g238 (n_226, wc28, n_180);
  not gc28 (wc28, n_183);
  or g239 (n_154, wc29, n_150);
  not gc29 (wc29, n_151);
  or g240 (n_227, wc30, n_185);
  not gc30 (wc30, n_188);
  or g241 (n_228, wc31, n_190);
  not gc31 (wc31, n_193);
  or g242 (n_159, wc32, n_155);
  not gc32 (wc32, n_156);
  or g243 (n_164, wc33, n_160);
  not gc33 (wc33, n_161);
  or g244 (n_169, wc34, n_165);
  not gc34 (wc34, n_166);
  or g245 (n_174, wc35, n_170);
  not gc35 (wc35, n_171);
  or g246 (n_179, wc36, n_175);
  not gc36 (wc36, n_176);
  or g247 (n_184, wc37, n_180);
  not gc37 (wc37, n_181);
  or g248 (n_189, wc38, n_185);
  not gc38 (wc38, n_186);
  or g249 (n_194, n_190, wc39);
  not gc39 (wc39, n_191);
  or g250 (n_199, n_195, wc40);
  not gc40 (wc40, n_196);
  or g251 (n_204, n_200, wc41);
  not gc41 (wc41, n_201);
  or g252 (n_209, n_205, wc42);
  not gc42 (wc42, n_206);
  or g253 (n_214, n_210, wc43);
  not gc43 (wc43, n_211);
endmodule

module csa_tree_add_104_26_group_173_GENERIC(in_0, in_1, in_2, out_0);
  input [8:0] in_0;
  input [1:0] in_1;
  input [15:0] in_2;
  output [15:0] out_0;
  wire [8:0] in_0;
  wire [1:0] in_1;
  wire [15:0] in_2;
  wire [15:0] out_0;
  csa_tree_add_104_26_group_173_GENERIC_REAL g1(.in_0 (in_0), .in_1
       (in_1), .in_2 (in_2), .out_0 (out_0));
endmodule

module csa_tree_add_116_28_group_175_GENERIC_REAL(in_0, in_1, in_2,
     out_0);
// synthesis_equation "assign out_0 = ( $signed(in_2) + ( $signed(in_0) * $signed(in_1) )  )  ;"
  input [15:0] in_0, in_2;
  input [1:0] in_1;
  output [15:0] out_0;
  wire [15:0] in_0, in_2;
  wire [1:0] in_1;
  wire [15:0] out_0;
  wire n_51, n_52, n_53, n_54, n_55, n_56, n_57, n_58;
  wire n_59, n_60, n_61, n_62, n_63, n_64, n_65, n_66;
  wire n_67, n_68, n_69, n_70, n_71, n_72, n_73, n_74;
  wire n_75, n_76, n_77, n_78, n_79, n_80, n_81, n_83;
  wire n_87, n_91, n_92, n_96, n_97, n_98, n_99, n_100;
  wire n_101, n_102, n_103, n_104, n_105, n_106, n_107, n_108;
  wire n_109, n_110, n_111, n_112, n_113, n_114, n_115, n_116;
  wire n_117, n_118, n_119, n_120, n_121, n_122, n_123, n_124;
  wire n_125, n_126, n_127, n_128, n_129, n_130, n_131, n_132;
  wire n_133, n_134, n_135, n_136, n_137, n_138, n_139, n_140;
  wire n_146, n_147, n_148, n_149, n_150, n_151, n_152, n_153;
  wire n_154, n_155, n_156, n_157, n_158, n_161, n_170, n_172;
  wire n_175, n_176, n_177, n_178, n_180, n_181, n_182, n_183;
  wire n_185, n_186, n_187, n_188, n_190, n_191, n_192, n_193;
  wire n_195, n_196, n_197, n_198, n_200, n_201, n_202, n_203;
  wire n_205, n_206, n_207, n_208, n_210, n_211, n_212, n_213;
  wire n_215, n_216, n_217, n_218, n_220, n_221, n_222, n_223;
  wire n_225, n_226, n_227, n_228, n_230, n_231, n_232, n_233;
  wire n_235, n_236, n_237, n_238, n_240, n_241, n_242, n_243;
  wire n_245, n_246, n_247, n_248, n_249, n_250, n_251, n_252;
  wire n_253, n_254, n_255, n_256, n_257, n_258, n_259, n_260;
  xor g3 (n_87, in_1[1], in_1[0]);
  xor g9 (n_91, in_1[1], in_0[0]);
  and g13 (n_66, in_0[0], in_1[0]);
  xor g14 (n_96, in_1[1], in_0[1]);
  nand g15 (n_97, n_96, in_1[0]);
  nand g16 (n_98, n_91, n_92);
  nand g17 (n_65, n_97, n_98);
  xor g18 (n_99, in_1[1], in_0[2]);
  nand g19 (n_100, n_99, in_1[0]);
  nand g20 (n_101, n_96, n_92);
  nand g21 (n_64, n_100, n_101);
  xor g22 (n_102, in_1[1], in_0[3]);
  nand g23 (n_103, n_102, in_1[0]);
  nand g24 (n_104, n_99, n_92);
  nand g25 (n_147, n_103, n_104);
  xor g26 (n_105, in_1[1], in_0[4]);
  nand g27 (n_106, n_105, in_1[0]);
  nand g28 (n_107, n_102, n_92);
  nand g29 (n_148, n_106, n_107);
  xor g30 (n_108, in_1[1], in_0[5]);
  nand g31 (n_109, n_108, in_1[0]);
  nand g32 (n_110, n_105, n_92);
  nand g33 (n_149, n_109, n_110);
  xor g34 (n_111, in_1[1], in_0[6]);
  nand g35 (n_112, n_111, in_1[0]);
  nand g36 (n_113, n_108, n_92);
  nand g37 (n_150, n_112, n_113);
  xor g38 (n_114, in_1[1], in_0[7]);
  nand g39 (n_115, n_114, in_1[0]);
  nand g40 (n_116, n_111, n_92);
  nand g41 (n_151, n_115, n_116);
  xor g42 (n_117, in_1[1], in_0[8]);
  nand g43 (n_118, n_117, in_1[0]);
  nand g44 (n_119, n_114, n_92);
  nand g45 (n_152, n_118, n_119);
  xor g46 (n_120, in_1[1], in_0[9]);
  nand g47 (n_121, n_120, in_1[0]);
  nand g48 (n_122, n_117, n_92);
  nand g49 (n_153, n_121, n_122);
  xor g50 (n_123, in_1[1], in_0[10]);
  nand g51 (n_124, n_123, in_1[0]);
  nand g52 (n_125, n_120, n_92);
  nand g53 (n_154, n_124, n_125);
  xor g54 (n_126, in_1[1], in_0[11]);
  nand g55 (n_127, n_126, in_1[0]);
  nand g56 (n_128, n_123, n_92);
  nand g57 (n_155, n_127, n_128);
  xor g58 (n_129, in_1[1], in_0[12]);
  nand g59 (n_130, n_129, in_1[0]);
  nand g60 (n_131, n_126, n_92);
  nand g61 (n_156, n_130, n_131);
  xor g62 (n_132, in_1[1], in_0[13]);
  nand g63 (n_133, n_132, in_1[0]);
  nand g64 (n_134, n_129, n_92);
  nand g65 (n_157, n_133, n_134);
  xor g66 (n_135, in_1[1], in_0[14]);
  nand g67 (n_136, n_135, in_1[0]);
  nand g68 (n_137, n_132, n_92);
  nand g69 (n_158, n_136, n_137);
  xor g70 (n_138, in_1[1], in_0[15]);
  nand g71 (n_139, n_138, in_1[0]);
  nand g72 (n_140, n_135, n_92);
  nand g73 (n_161, n_139, n_140);
  xor g93 (n_81, in_2[1], n_83);
  and g94 (n_146, in_2[1], n_83);
  xor g95 (n_80, in_2[2], n_146);
  and g96 (n_63, in_2[2], n_146);
  xor g97 (n_79, in_2[3], n_147);
  and g98 (n_62, in_2[3], n_147);
  xor g99 (n_78, in_2[4], n_148);
  and g100 (n_61, in_2[4], n_148);
  xor g101 (n_77, in_2[5], n_149);
  and g102 (n_60, in_2[5], n_149);
  xor g103 (n_76, in_2[6], n_150);
  and g104 (n_59, in_2[6], n_150);
  xor g105 (n_75, in_2[7], n_151);
  and g106 (n_58, in_2[7], n_151);
  xor g107 (n_74, in_2[8], n_152);
  and g108 (n_57, in_2[8], n_152);
  xor g109 (n_73, in_2[9], n_153);
  and g110 (n_56, in_2[9], n_153);
  xor g111 (n_72, in_2[10], n_154);
  and g112 (n_55, in_2[10], n_154);
  xor g113 (n_71, in_2[11], n_155);
  and g114 (n_54, in_2[11], n_155);
  xor g115 (n_70, in_2[12], n_156);
  and g116 (n_53, in_2[12], n_156);
  xor g117 (n_69, in_2[13], n_157);
  and g118 (n_52, in_2[13], n_157);
  xor g119 (n_68, in_2[14], n_158);
  and g120 (n_51, in_2[14], n_158);
  xor g122 (n_67, in_2[15], n_161);
  nand g131 (n_170, n_66, in_2[0]);
  nor g134 (n_172, n_65, n_81);
  nand g135 (n_175, n_65, n_81);
  nor g136 (n_177, n_64, n_80);
  nand g137 (n_180, n_64, n_80);
  nor g138 (n_182, n_63, n_79);
  nand g139 (n_185, n_63, n_79);
  nor g140 (n_187, n_62, n_78);
  nand g141 (n_190, n_62, n_78);
  nor g142 (n_192, n_61, n_77);
  nand g143 (n_195, n_61, n_77);
  nor g144 (n_197, n_60, n_76);
  nand g145 (n_200, n_60, n_76);
  nor g146 (n_202, n_59, n_75);
  nand g147 (n_205, n_59, n_75);
  nor g148 (n_207, n_58, n_74);
  nand g149 (n_210, n_58, n_74);
  nor g150 (n_212, n_57, n_73);
  nand g151 (n_215, n_57, n_73);
  nor g152 (n_217, n_56, n_72);
  nand g153 (n_220, n_56, n_72);
  nor g154 (n_222, n_55, n_71);
  nand g155 (n_225, n_55, n_71);
  nor g156 (n_227, n_54, n_70);
  nand g157 (n_230, n_54, n_70);
  nor g158 (n_232, n_53, n_69);
  nand g159 (n_235, n_53, n_69);
  nor g160 (n_237, n_52, n_68);
  nand g161 (n_240, n_52, n_68);
  nand g166 (n_178, n_175, n_176);
  nand g169 (n_183, n_180, n_181);
  nand g172 (n_188, n_185, n_186);
  nand g175 (n_193, n_190, n_191);
  nand g178 (n_198, n_195, n_196);
  nand g181 (n_203, n_200, n_201);
  nand g184 (n_208, n_205, n_206);
  nand g187 (n_213, n_210, n_211);
  nand g190 (n_218, n_215, n_216);
  nand g193 (n_223, n_220, n_221);
  nand g196 (n_228, n_225, n_226);
  nand g199 (n_233, n_230, n_231);
  nand g202 (n_238, n_235, n_236);
  nand g80 (n_243, n_240, n_241);
  xnor g87 (out_0[2], n_178, n_247);
  xnor g89 (out_0[3], n_183, n_248);
  xnor g91 (out_0[4], n_188, n_249);
  xnor g203 (out_0[5], n_193, n_250);
  xnor g205 (out_0[6], n_198, n_251);
  xnor g207 (out_0[7], n_203, n_252);
  xnor g209 (out_0[8], n_208, n_253);
  xnor g211 (out_0[9], n_213, n_254);
  xnor g213 (out_0[10], n_218, n_255);
  xnor g215 (out_0[11], n_223, n_256);
  xnor g217 (out_0[12], n_228, n_257);
  xnor g219 (out_0[13], n_233, n_258);
  xnor g221 (out_0[14], n_238, n_259);
  xnor g223 (out_0[15], n_243, n_260);
  xor g224 (out_0[0], in_2[0], n_66);
  and g226 (n_92, wc, n_87);
  not gc (wc, in_1[0]);
  and g228 (n_83, in_1[1], wc0);
  not gc0 (wc0, n_66);
  and g230 (n_242, n_51, n_67);
  or g231 (n_245, n_51, n_67);
  or g232 (n_176, n_170, n_172);
  or g233 (n_246, wc1, n_172);
  not gc1 (wc1, n_175);
  xor g234 (out_0[1], n_170, n_246);
  or g235 (n_247, wc2, n_177);
  not gc2 (wc2, n_180);
  or g236 (n_248, wc3, n_182);
  not gc3 (wc3, n_185);
  or g237 (n_249, wc4, n_187);
  not gc4 (wc4, n_190);
  or g238 (n_250, wc5, n_192);
  not gc5 (wc5, n_195);
  or g239 (n_251, wc6, n_197);
  not gc6 (wc6, n_200);
  or g240 (n_252, wc7, n_202);
  not gc7 (wc7, n_205);
  or g241 (n_253, wc8, n_207);
  not gc8 (wc8, n_210);
  or g242 (n_254, wc9, n_212);
  not gc9 (wc9, n_215);
  or g243 (n_255, wc10, n_217);
  not gc10 (wc10, n_220);
  or g244 (n_256, wc11, n_222);
  not gc11 (wc11, n_225);
  or g245 (n_257, wc12, n_227);
  not gc12 (wc12, n_230);
  or g246 (n_258, wc13, n_232);
  not gc13 (wc13, n_235);
  or g247 (n_259, wc14, n_237);
  not gc14 (wc14, n_240);
  or g248 (n_181, wc15, n_177);
  not gc15 (wc15, n_178);
  or g249 (n_260, wc16, n_242);
  not gc16 (wc16, n_245);
  or g250 (n_186, wc17, n_182);
  not gc17 (wc17, n_183);
  or g251 (n_191, wc18, n_187);
  not gc18 (wc18, n_188);
  or g252 (n_196, wc19, n_192);
  not gc19 (wc19, n_193);
  or g253 (n_201, wc20, n_197);
  not gc20 (wc20, n_198);
  or g254 (n_206, wc21, n_202);
  not gc21 (wc21, n_203);
  or g255 (n_211, wc22, n_207);
  not gc22 (wc22, n_208);
  or g256 (n_216, wc23, n_212);
  not gc23 (wc23, n_213);
  or g257 (n_221, wc24, n_217);
  not gc24 (wc24, n_218);
  or g258 (n_226, wc25, n_222);
  not gc25 (wc25, n_223);
  or g259 (n_231, wc26, n_227);
  not gc26 (wc26, n_228);
  or g260 (n_236, wc27, n_232);
  not gc27 (wc27, n_233);
  or g261 (n_241, wc28, n_237);
  not gc28 (wc28, n_238);
endmodule

module csa_tree_add_116_28_group_175_GENERIC(in_0, in_1, in_2, out_0);
  input [15:0] in_0, in_2;
  input [1:0] in_1;
  output [15:0] out_0;
  wire [15:0] in_0, in_2;
  wire [1:0] in_1;
  wire [15:0] out_0;
  csa_tree_add_116_28_group_175_GENERIC_REAL g1(.in_0 (in_0), .in_1
       (in_1), .in_2 (in_2), .out_0 (out_0));
endmodule

