module csa_tree_add_38_13_group_93_GENERIC_REAL(in_0, in_1, in_2,
     out_0);
// synthesis_equation "assign out_0 = ( $signed(in_2) + ( $signed(in_0) * $signed(in_1) )  )  ;"
  input [1:0] in_0;
  input [8:0] in_1;
  input [11:0] in_2;
  output [11:0] out_0;
  wire [1:0] in_0;
  wire [8:0] in_1;
  wire [11:0] in_2;
  wire [11:0] out_0;
  wire n_38, n_39, n_40, n_41, n_42, n_43, n_44, n_45;
  wire n_46, n_47, n_49, n_50, n_51, n_52, n_53, n_54;
  wire n_55, n_56, n_57, n_58, n_60, n_64, n_68, n_69;
  wire n_73, n_74, n_75, n_76, n_77, n_78, n_79, n_80;
  wire n_81, n_82, n_83, n_84, n_85, n_86, n_87, n_88;
  wire n_89, n_90, n_91, n_92, n_93, n_94, n_95, n_96;
  wire n_99, n_100, n_106, n_107, n_108, n_109, n_110, n_111;
  wire n_112, n_113, n_120, n_124, n_126, n_129, n_130, n_131;
  wire n_132, n_134, n_135, n_136, n_137, n_139, n_140, n_141;
  wire n_143, n_144, n_145, n_146, n_148, n_149, n_150, n_151;
  wire n_153, n_154, n_155, n_156, n_158, n_159, n_160, n_161;
  wire n_163, n_164, n_165, n_166, n_168, n_169, n_170, n_171;
  wire n_173, n_174, n_175, n_176, n_178, n_179, n_180, n_181;
  wire n_182, n_183, n_184, n_185, n_186, n_187, n_188, n_189;
  xor g3 (n_64, in_0[1], in_0[0]);
  xor g9 (n_68, in_0[1], in_1[0]);
  and g13 (n_47, in_1[0], in_0[0]);
  xor g14 (n_73, in_0[1], in_1[1]);
  nand g15 (n_74, n_73, in_0[0]);
  nand g16 (n_75, n_68, n_69);
  nand g17 (n_46, n_74, n_75);
  xor g18 (n_76, in_0[1], in_1[2]);
  nand g19 (n_77, n_76, in_0[0]);
  nand g20 (n_78, n_73, n_69);
  nand g21 (n_45, n_77, n_78);
  xor g22 (n_79, in_0[1], in_1[3]);
  nand g23 (n_80, n_79, in_0[0]);
  nand g24 (n_81, n_76, n_69);
  nand g25 (n_108, n_80, n_81);
  xor g26 (n_82, in_0[1], in_1[4]);
  nand g27 (n_83, n_82, in_0[0]);
  nand g28 (n_84, n_79, n_69);
  nand g29 (n_109, n_83, n_84);
  xor g30 (n_85, in_0[1], in_1[5]);
  nand g31 (n_86, n_85, in_0[0]);
  nand g32 (n_87, n_82, n_69);
  nand g33 (n_110, n_86, n_87);
  xor g34 (n_88, in_0[1], in_1[6]);
  nand g35 (n_89, n_88, in_0[0]);
  nand g36 (n_90, n_85, n_69);
  nand g37 (n_111, n_89, n_90);
  xor g38 (n_91, in_0[1], in_1[7]);
  nand g39 (n_92, n_91, in_0[0]);
  nand g40 (n_93, n_88, n_69);
  nand g41 (n_112, n_92, n_93);
  xor g42 (n_94, in_0[1], in_1[8]);
  nand g43 (n_95, n_94, in_0[0]);
  nand g44 (n_96, n_91, n_69);
  nand g45 (n_113, n_95, n_96);
  nand g48 (n_99, n_94, n_69);
  nand g49 (n_100, n_95, n_99);
  xor g65 (n_58, in_2[1], n_106);
  and g66 (n_107, in_2[1], n_106);
  xor g67 (n_57, in_2[2], n_107);
  and g68 (n_44, in_2[2], n_107);
  xor g69 (n_56, in_2[3], n_108);
  and g70 (n_43, in_2[3], n_108);
  xor g71 (n_55, in_2[4], n_109);
  and g72 (n_42, in_2[4], n_109);
  xor g73 (n_54, in_2[5], n_110);
  and g74 (n_41, in_2[5], n_110);
  xor g75 (n_53, in_2[6], n_111);
  and g76 (n_40, in_2[6], n_111);
  xor g77 (n_52, in_2[7], n_112);
  and g78 (n_39, in_2[7], n_112);
  xor g79 (n_51, in_2[8], n_113);
  and g80 (n_38, in_2[8], n_113);
  nand g93 (n_124, n_47, in_2[0]);
  nor g96 (n_126, n_46, n_58);
  nand g97 (n_129, n_46, n_58);
  nor g98 (n_131, n_45, n_57);
  nand g99 (n_134, n_45, n_57);
  nor g100 (n_136, n_44, n_56);
  nand g101 (n_139, n_44, n_56);
  nor g102 (n_60, n_43, n_55);
  nand g103 (n_143, n_43, n_55);
  nor g104 (n_145, n_42, n_54);
  nand g105 (n_148, n_42, n_54);
  nor g106 (n_150, n_41, n_53);
  nand g107 (n_153, n_41, n_53);
  nor g108 (n_155, n_40, n_52);
  nand g109 (n_158, n_40, n_52);
  nor g110 (n_160, n_39, n_51);
  nand g111 (n_163, n_39, n_51);
  nor g112 (n_165, n_38, n_50);
  nand g113 (n_168, n_38, n_50);
  nand g120 (n_132, n_129, n_130);
  nand g123 (n_137, n_134, n_135);
  nand g126 (n_141, n_139, n_140);
  nand g129 (n_146, n_143, n_144);
  nand g132 (n_151, n_148, n_149);
  nand g135 (n_156, n_153, n_154);
  nand g138 (n_161, n_158, n_159);
  nand g141 (n_166, n_163, n_164);
  nand g57 (n_171, n_168, n_169);
  nand g60 (n_176, n_173, n_174);
  xnor g144 (out_0[2], n_132, n_180);
  xnor g146 (out_0[3], n_137, n_181);
  xnor g148 (out_0[4], n_141, n_182);
  xnor g150 (out_0[5], n_146, n_183);
  xnor g152 (out_0[6], n_151, n_184);
  xnor g154 (out_0[7], n_156, n_185);
  xnor g156 (out_0[8], n_161, n_186);
  xnor g158 (out_0[9], n_166, n_187);
  xnor g160 (out_0[10], n_171, n_188);
  xnor g162 (out_0[11], n_176, n_189);
  xor g163 (out_0[0], in_2[0], n_47);
  and g167 (n_69, wc, n_64);
  not gc (wc, in_0[0]);
  and g169 (n_175, in_2[10], wc0);
  not gc0 (wc0, in_2[11]);
  or g170 (n_178, in_2[10], wc1);
  not gc1 (wc1, in_2[11]);
  and g171 (n_106, in_0[1], wc2);
  not gc2 (wc2, n_47);
  or g173 (n_189, wc3, n_175);
  not gc3 (wc3, n_178);
  xor g174 (n_50, n_100, in_2[9]);
  or g175 (n_120, wc4, n_100);
  not gc4 (wc4, in_2[9]);
  or g176 (n_49, in_2[9], wc5, wc6);
  not gc6 (wc6, n_100);
  not gc5 (wc5, n_120);
  or g177 (n_130, n_124, n_126);
  or g178 (n_179, wc7, n_126);
  not gc7 (wc7, n_129);
  and g179 (n_170, in_2[10], wc8);
  not gc8 (wc8, n_49);
  or g180 (n_173, in_2[10], wc9);
  not gc9 (wc9, n_49);
  xor g181 (out_0[1], n_124, n_179);
  or g182 (n_180, wc10, n_131);
  not gc10 (wc10, n_134);
  or g183 (n_181, wc11, n_136);
  not gc11 (wc11, n_139);
  or g184 (n_182, wc12, n_60);
  not gc12 (wc12, n_143);
  or g185 (n_183, wc13, n_145);
  not gc13 (wc13, n_148);
  or g186 (n_184, wc14, n_150);
  not gc14 (wc14, n_153);
  or g187 (n_185, wc15, n_155);
  not gc15 (wc15, n_158);
  or g188 (n_186, wc16, n_160);
  not gc16 (wc16, n_163);
  or g189 (n_135, wc17, n_131);
  not gc17 (wc17, n_132);
  or g190 (n_187, wc18, n_165);
  not gc18 (wc18, n_168);
  or g191 (n_188, wc19, n_170);
  not gc19 (wc19, n_173);
  or g192 (n_140, wc20, n_136);
  not gc20 (wc20, n_137);
  or g193 (n_144, wc21, n_60);
  not gc21 (wc21, n_141);
  or g194 (n_149, wc22, n_145);
  not gc22 (wc22, n_146);
  or g195 (n_154, wc23, n_150);
  not gc23 (wc23, n_151);
  or g196 (n_159, wc24, n_155);
  not gc24 (wc24, n_156);
  or g197 (n_164, wc25, n_160);
  not gc25 (wc25, n_161);
  or g198 (n_169, wc26, n_165);
  not gc26 (wc26, n_166);
  or g199 (n_174, n_170, wc27);
  not gc27 (wc27, n_171);
endmodule

module csa_tree_add_38_13_group_93_GENERIC(in_0, in_1, in_2, out_0);
  input [1:0] in_0;
  input [8:0] in_1;
  input [11:0] in_2;
  output [11:0] out_0;
  wire [1:0] in_0;
  wire [8:0] in_1;
  wire [11:0] in_2;
  wire [11:0] out_0;
  csa_tree_add_38_13_group_93_GENERIC_REAL g1(.in_0 (in_0), .in_1
       (in_1), .in_2 (in_2), .out_0 (out_0));
endmodule

module csa_tree_add_38_13_group_93_154_GENERIC_REAL(in_0, in_1, in_2,
     out_0);
// synthesis_equation "assign out_0 = ( $signed(in_2) + ( $signed(in_0) * $signed(in_1) )  )  ;"
  input [1:0] in_0;
  input [8:0] in_1;
  input [11:0] in_2;
  output [11:0] out_0;
  wire [1:0] in_0;
  wire [8:0] in_1;
  wire [11:0] in_2;
  wire [11:0] out_0;
  wire n_38, n_39, n_40, n_41, n_42, n_43, n_44, n_45;
  wire n_46, n_47, n_49, n_50, n_51, n_52, n_53, n_54;
  wire n_55, n_56, n_57, n_58, n_60, n_64, n_68, n_69;
  wire n_73, n_74, n_75, n_76, n_77, n_78, n_79, n_80;
  wire n_81, n_82, n_83, n_84, n_85, n_86, n_87, n_88;
  wire n_89, n_90, n_91, n_92, n_93, n_94, n_95, n_96;
  wire n_99, n_100, n_106, n_107, n_108, n_109, n_110, n_111;
  wire n_112, n_113, n_120, n_124, n_126, n_129, n_130, n_131;
  wire n_132, n_134, n_135, n_136, n_137, n_139, n_140, n_141;
  wire n_143, n_144, n_145, n_146, n_148, n_149, n_150, n_151;
  wire n_153, n_154, n_155, n_156, n_158, n_159, n_160, n_161;
  wire n_163, n_164, n_165, n_166, n_168, n_169, n_170, n_171;
  wire n_173, n_174, n_175, n_176, n_178, n_179, n_180, n_181;
  wire n_182, n_183, n_184, n_185, n_186, n_187, n_188, n_189;
  xor g3 (n_64, in_0[1], in_0[0]);
  xor g9 (n_68, in_0[1], in_1[0]);
  and g13 (n_47, in_1[0], in_0[0]);
  xor g14 (n_73, in_0[1], in_1[1]);
  nand g15 (n_74, n_73, in_0[0]);
  nand g16 (n_75, n_68, n_69);
  nand g17 (n_46, n_74, n_75);
  xor g18 (n_76, in_0[1], in_1[2]);
  nand g19 (n_77, n_76, in_0[0]);
  nand g20 (n_78, n_73, n_69);
  nand g21 (n_45, n_77, n_78);
  xor g22 (n_79, in_0[1], in_1[3]);
  nand g23 (n_80, n_79, in_0[0]);
  nand g24 (n_81, n_76, n_69);
  nand g25 (n_108, n_80, n_81);
  xor g26 (n_82, in_0[1], in_1[4]);
  nand g27 (n_83, n_82, in_0[0]);
  nand g28 (n_84, n_79, n_69);
  nand g29 (n_109, n_83, n_84);
  xor g30 (n_85, in_0[1], in_1[5]);
  nand g31 (n_86, n_85, in_0[0]);
  nand g32 (n_87, n_82, n_69);
  nand g33 (n_110, n_86, n_87);
  xor g34 (n_88, in_0[1], in_1[6]);
  nand g35 (n_89, n_88, in_0[0]);
  nand g36 (n_90, n_85, n_69);
  nand g37 (n_111, n_89, n_90);
  xor g38 (n_91, in_0[1], in_1[7]);
  nand g39 (n_92, n_91, in_0[0]);
  nand g40 (n_93, n_88, n_69);
  nand g41 (n_112, n_92, n_93);
  xor g42 (n_94, in_0[1], in_1[8]);
  nand g43 (n_95, n_94, in_0[0]);
  nand g44 (n_96, n_91, n_69);
  nand g45 (n_113, n_95, n_96);
  nand g48 (n_99, n_94, n_69);
  nand g49 (n_100, n_95, n_99);
  xor g65 (n_58, in_2[1], n_106);
  and g66 (n_107, in_2[1], n_106);
  xor g67 (n_57, in_2[2], n_107);
  and g68 (n_44, in_2[2], n_107);
  xor g69 (n_56, in_2[3], n_108);
  and g70 (n_43, in_2[3], n_108);
  xor g71 (n_55, in_2[4], n_109);
  and g72 (n_42, in_2[4], n_109);
  xor g73 (n_54, in_2[5], n_110);
  and g74 (n_41, in_2[5], n_110);
  xor g75 (n_53, in_2[6], n_111);
  and g76 (n_40, in_2[6], n_111);
  xor g77 (n_52, in_2[7], n_112);
  and g78 (n_39, in_2[7], n_112);
  xor g79 (n_51, in_2[8], n_113);
  and g80 (n_38, in_2[8], n_113);
  nand g93 (n_124, n_47, in_2[0]);
  nor g96 (n_126, n_46, n_58);
  nand g97 (n_129, n_46, n_58);
  nor g98 (n_131, n_45, n_57);
  nand g99 (n_134, n_45, n_57);
  nor g100 (n_136, n_44, n_56);
  nand g101 (n_139, n_44, n_56);
  nor g102 (n_60, n_43, n_55);
  nand g103 (n_143, n_43, n_55);
  nor g104 (n_145, n_42, n_54);
  nand g105 (n_148, n_42, n_54);
  nor g106 (n_150, n_41, n_53);
  nand g107 (n_153, n_41, n_53);
  nor g108 (n_155, n_40, n_52);
  nand g109 (n_158, n_40, n_52);
  nor g110 (n_160, n_39, n_51);
  nand g111 (n_163, n_39, n_51);
  nor g112 (n_165, n_38, n_50);
  nand g113 (n_168, n_38, n_50);
  nand g120 (n_132, n_129, n_130);
  nand g123 (n_137, n_134, n_135);
  nand g126 (n_141, n_139, n_140);
  nand g129 (n_146, n_143, n_144);
  nand g132 (n_151, n_148, n_149);
  nand g135 (n_156, n_153, n_154);
  nand g138 (n_161, n_158, n_159);
  nand g141 (n_166, n_163, n_164);
  nand g57 (n_171, n_168, n_169);
  nand g60 (n_176, n_173, n_174);
  xnor g144 (out_0[2], n_132, n_180);
  xnor g146 (out_0[3], n_137, n_181);
  xnor g148 (out_0[4], n_141, n_182);
  xnor g150 (out_0[5], n_146, n_183);
  xnor g152 (out_0[6], n_151, n_184);
  xnor g154 (out_0[7], n_156, n_185);
  xnor g156 (out_0[8], n_161, n_186);
  xnor g158 (out_0[9], n_166, n_187);
  xnor g160 (out_0[10], n_171, n_188);
  xnor g162 (out_0[11], n_176, n_189);
  xor g163 (out_0[0], in_2[0], n_47);
  and g167 (n_69, wc, n_64);
  not gc (wc, in_0[0]);
  and g169 (n_175, in_2[10], wc0);
  not gc0 (wc0, in_2[11]);
  or g170 (n_178, in_2[10], wc1);
  not gc1 (wc1, in_2[11]);
  and g171 (n_106, in_0[1], wc2);
  not gc2 (wc2, n_47);
  or g173 (n_189, wc3, n_175);
  not gc3 (wc3, n_178);
  xor g174 (n_50, n_100, in_2[9]);
  or g175 (n_120, wc4, n_100);
  not gc4 (wc4, in_2[9]);
  or g176 (n_49, in_2[9], wc5, wc6);
  not gc6 (wc6, n_100);
  not gc5 (wc5, n_120);
  or g177 (n_130, n_124, n_126);
  or g178 (n_179, wc7, n_126);
  not gc7 (wc7, n_129);
  and g179 (n_170, in_2[10], wc8);
  not gc8 (wc8, n_49);
  or g180 (n_173, in_2[10], wc9);
  not gc9 (wc9, n_49);
  xor g181 (out_0[1], n_124, n_179);
  or g182 (n_180, wc10, n_131);
  not gc10 (wc10, n_134);
  or g183 (n_181, wc11, n_136);
  not gc11 (wc11, n_139);
  or g184 (n_182, wc12, n_60);
  not gc12 (wc12, n_143);
  or g185 (n_183, wc13, n_145);
  not gc13 (wc13, n_148);
  or g186 (n_184, wc14, n_150);
  not gc14 (wc14, n_153);
  or g187 (n_185, wc15, n_155);
  not gc15 (wc15, n_158);
  or g188 (n_186, wc16, n_160);
  not gc16 (wc16, n_163);
  or g189 (n_135, wc17, n_131);
  not gc17 (wc17, n_132);
  or g190 (n_187, wc18, n_165);
  not gc18 (wc18, n_168);
  or g191 (n_188, wc19, n_170);
  not gc19 (wc19, n_173);
  or g192 (n_140, wc20, n_136);
  not gc20 (wc20, n_137);
  or g193 (n_144, wc21, n_60);
  not gc21 (wc21, n_141);
  or g194 (n_149, wc22, n_145);
  not gc22 (wc22, n_146);
  or g195 (n_154, wc23, n_150);
  not gc23 (wc23, n_151);
  or g196 (n_159, wc24, n_155);
  not gc24 (wc24, n_156);
  or g197 (n_164, wc25, n_160);
  not gc25 (wc25, n_161);
  or g198 (n_169, wc26, n_165);
  not gc26 (wc26, n_166);
  or g199 (n_174, n_170, wc27);
  not gc27 (wc27, n_171);
endmodule

module csa_tree_add_38_13_group_93_154_GENERIC(in_0, in_1, in_2, out_0);
  input [1:0] in_0;
  input [8:0] in_1;
  input [11:0] in_2;
  output [11:0] out_0;
  wire [1:0] in_0;
  wire [8:0] in_1;
  wire [11:0] in_2;
  wire [11:0] out_0;
  csa_tree_add_38_13_group_93_154_GENERIC_REAL g1(.in_0 (in_0), .in_1
       (in_1), .in_2 (in_2), .out_0 (out_0));
endmodule

module csa_tree_add_38_13_group_93_155_GENERIC_REAL(in_0, in_1, in_2,
     out_0);
// synthesis_equation "assign out_0 = ( $signed(in_2) + ( $signed(in_0) * $signed(in_1) )  )  ;"
  input [1:0] in_0;
  input [8:0] in_1;
  input [11:0] in_2;
  output [11:0] out_0;
  wire [1:0] in_0;
  wire [8:0] in_1;
  wire [11:0] in_2;
  wire [11:0] out_0;
  wire n_38, n_39, n_40, n_41, n_42, n_43, n_44, n_45;
  wire n_46, n_47, n_49, n_50, n_51, n_52, n_53, n_54;
  wire n_55, n_56, n_57, n_58, n_60, n_64, n_68, n_69;
  wire n_73, n_74, n_75, n_76, n_77, n_78, n_79, n_80;
  wire n_81, n_82, n_83, n_84, n_85, n_86, n_87, n_88;
  wire n_89, n_90, n_91, n_92, n_93, n_94, n_95, n_96;
  wire n_99, n_100, n_106, n_107, n_108, n_109, n_110, n_111;
  wire n_112, n_113, n_120, n_124, n_126, n_129, n_130, n_131;
  wire n_132, n_134, n_135, n_136, n_137, n_139, n_140, n_141;
  wire n_143, n_144, n_145, n_146, n_148, n_149, n_150, n_151;
  wire n_153, n_154, n_155, n_156, n_158, n_159, n_160, n_161;
  wire n_163, n_164, n_165, n_166, n_168, n_169, n_170, n_171;
  wire n_173, n_174, n_175, n_176, n_178, n_179, n_180, n_181;
  wire n_182, n_183, n_184, n_185, n_186, n_187, n_188, n_189;
  xor g3 (n_64, in_0[1], in_0[0]);
  xor g9 (n_68, in_0[1], in_1[0]);
  and g13 (n_47, in_1[0], in_0[0]);
  xor g14 (n_73, in_0[1], in_1[1]);
  nand g15 (n_74, n_73, in_0[0]);
  nand g16 (n_75, n_68, n_69);
  nand g17 (n_46, n_74, n_75);
  xor g18 (n_76, in_0[1], in_1[2]);
  nand g19 (n_77, n_76, in_0[0]);
  nand g20 (n_78, n_73, n_69);
  nand g21 (n_45, n_77, n_78);
  xor g22 (n_79, in_0[1], in_1[3]);
  nand g23 (n_80, n_79, in_0[0]);
  nand g24 (n_81, n_76, n_69);
  nand g25 (n_108, n_80, n_81);
  xor g26 (n_82, in_0[1], in_1[4]);
  nand g27 (n_83, n_82, in_0[0]);
  nand g28 (n_84, n_79, n_69);
  nand g29 (n_109, n_83, n_84);
  xor g30 (n_85, in_0[1], in_1[5]);
  nand g31 (n_86, n_85, in_0[0]);
  nand g32 (n_87, n_82, n_69);
  nand g33 (n_110, n_86, n_87);
  xor g34 (n_88, in_0[1], in_1[6]);
  nand g35 (n_89, n_88, in_0[0]);
  nand g36 (n_90, n_85, n_69);
  nand g37 (n_111, n_89, n_90);
  xor g38 (n_91, in_0[1], in_1[7]);
  nand g39 (n_92, n_91, in_0[0]);
  nand g40 (n_93, n_88, n_69);
  nand g41 (n_112, n_92, n_93);
  xor g42 (n_94, in_0[1], in_1[8]);
  nand g43 (n_95, n_94, in_0[0]);
  nand g44 (n_96, n_91, n_69);
  nand g45 (n_113, n_95, n_96);
  nand g48 (n_99, n_94, n_69);
  nand g49 (n_100, n_95, n_99);
  xor g65 (n_58, in_2[1], n_106);
  and g66 (n_107, in_2[1], n_106);
  xor g67 (n_57, in_2[2], n_107);
  and g68 (n_44, in_2[2], n_107);
  xor g69 (n_56, in_2[3], n_108);
  and g70 (n_43, in_2[3], n_108);
  xor g71 (n_55, in_2[4], n_109);
  and g72 (n_42, in_2[4], n_109);
  xor g73 (n_54, in_2[5], n_110);
  and g74 (n_41, in_2[5], n_110);
  xor g75 (n_53, in_2[6], n_111);
  and g76 (n_40, in_2[6], n_111);
  xor g77 (n_52, in_2[7], n_112);
  and g78 (n_39, in_2[7], n_112);
  xor g79 (n_51, in_2[8], n_113);
  and g80 (n_38, in_2[8], n_113);
  nand g93 (n_124, n_47, in_2[0]);
  nor g96 (n_126, n_46, n_58);
  nand g97 (n_129, n_46, n_58);
  nor g98 (n_131, n_45, n_57);
  nand g99 (n_134, n_45, n_57);
  nor g100 (n_136, n_44, n_56);
  nand g101 (n_139, n_44, n_56);
  nor g102 (n_60, n_43, n_55);
  nand g103 (n_143, n_43, n_55);
  nor g104 (n_145, n_42, n_54);
  nand g105 (n_148, n_42, n_54);
  nor g106 (n_150, n_41, n_53);
  nand g107 (n_153, n_41, n_53);
  nor g108 (n_155, n_40, n_52);
  nand g109 (n_158, n_40, n_52);
  nor g110 (n_160, n_39, n_51);
  nand g111 (n_163, n_39, n_51);
  nor g112 (n_165, n_38, n_50);
  nand g113 (n_168, n_38, n_50);
  nand g120 (n_132, n_129, n_130);
  nand g123 (n_137, n_134, n_135);
  nand g126 (n_141, n_139, n_140);
  nand g129 (n_146, n_143, n_144);
  nand g132 (n_151, n_148, n_149);
  nand g135 (n_156, n_153, n_154);
  nand g138 (n_161, n_158, n_159);
  nand g141 (n_166, n_163, n_164);
  nand g57 (n_171, n_168, n_169);
  nand g60 (n_176, n_173, n_174);
  xnor g144 (out_0[2], n_132, n_180);
  xnor g146 (out_0[3], n_137, n_181);
  xnor g148 (out_0[4], n_141, n_182);
  xnor g150 (out_0[5], n_146, n_183);
  xnor g152 (out_0[6], n_151, n_184);
  xnor g154 (out_0[7], n_156, n_185);
  xnor g156 (out_0[8], n_161, n_186);
  xnor g158 (out_0[9], n_166, n_187);
  xnor g160 (out_0[10], n_171, n_188);
  xnor g162 (out_0[11], n_176, n_189);
  xor g163 (out_0[0], in_2[0], n_47);
  and g167 (n_69, wc, n_64);
  not gc (wc, in_0[0]);
  and g169 (n_175, in_2[10], wc0);
  not gc0 (wc0, in_2[11]);
  or g170 (n_178, in_2[10], wc1);
  not gc1 (wc1, in_2[11]);
  and g171 (n_106, in_0[1], wc2);
  not gc2 (wc2, n_47);
  or g173 (n_189, wc3, n_175);
  not gc3 (wc3, n_178);
  xor g174 (n_50, n_100, in_2[9]);
  or g175 (n_120, wc4, n_100);
  not gc4 (wc4, in_2[9]);
  or g176 (n_49, in_2[9], wc5, wc6);
  not gc6 (wc6, n_100);
  not gc5 (wc5, n_120);
  or g177 (n_130, n_124, n_126);
  or g178 (n_179, wc7, n_126);
  not gc7 (wc7, n_129);
  and g179 (n_170, in_2[10], wc8);
  not gc8 (wc8, n_49);
  or g180 (n_173, in_2[10], wc9);
  not gc9 (wc9, n_49);
  xor g181 (out_0[1], n_124, n_179);
  or g182 (n_180, wc10, n_131);
  not gc10 (wc10, n_134);
  or g183 (n_181, wc11, n_136);
  not gc11 (wc11, n_139);
  or g184 (n_182, wc12, n_60);
  not gc12 (wc12, n_143);
  or g185 (n_183, wc13, n_145);
  not gc13 (wc13, n_148);
  or g186 (n_184, wc14, n_150);
  not gc14 (wc14, n_153);
  or g187 (n_185, wc15, n_155);
  not gc15 (wc15, n_158);
  or g188 (n_186, wc16, n_160);
  not gc16 (wc16, n_163);
  or g189 (n_135, wc17, n_131);
  not gc17 (wc17, n_132);
  or g190 (n_187, wc18, n_165);
  not gc18 (wc18, n_168);
  or g191 (n_188, wc19, n_170);
  not gc19 (wc19, n_173);
  or g192 (n_140, wc20, n_136);
  not gc20 (wc20, n_137);
  or g193 (n_144, wc21, n_60);
  not gc21 (wc21, n_141);
  or g194 (n_149, wc22, n_145);
  not gc22 (wc22, n_146);
  or g195 (n_154, wc23, n_150);
  not gc23 (wc23, n_151);
  or g196 (n_159, wc24, n_155);
  not gc24 (wc24, n_156);
  or g197 (n_164, wc25, n_160);
  not gc25 (wc25, n_161);
  or g198 (n_169, wc26, n_165);
  not gc26 (wc26, n_166);
  or g199 (n_174, n_170, wc27);
  not gc27 (wc27, n_171);
endmodule

module csa_tree_add_38_13_group_93_155_GENERIC(in_0, in_1, in_2, out_0);
  input [1:0] in_0;
  input [8:0] in_1;
  input [11:0] in_2;
  output [11:0] out_0;
  wire [1:0] in_0;
  wire [8:0] in_1;
  wire [11:0] in_2;
  wire [11:0] out_0;
  csa_tree_add_38_13_group_93_155_GENERIC_REAL g1(.in_0 (in_0), .in_1
       (in_1), .in_2 (in_2), .out_0 (out_0));
endmodule

module csa_tree_add_52_27_group_97_GENERIC_REAL(in_0, in_1, in_2,
     out_0);
// synthesis_equation "assign out_0 = ( ( $signed(in_1) + $signed(in_2) )  + $signed(in_0) )  ;"
  input [10:0] in_0, in_1, in_2;
  output [10:0] out_0;
  wire [10:0] in_0, in_1, in_2;
  wire [10:0] out_0;
  wire n_45, n_46, n_47, n_48, n_49, n_50, n_51, n_52;
  wire n_53, n_55, n_56, n_57, n_58, n_59, n_60, n_61;
  wire n_62, n_63, n_64, n_65, n_66, n_67, n_72, n_73;
  wire n_74, n_75, n_76, n_77, n_78, n_79, n_80, n_81;
  wire n_82, n_83, n_84, n_85, n_86, n_87, n_88, n_89;
  wire n_90, n_91, n_92, n_93, n_94, n_95, n_96, n_97;
  wire n_98, n_99, n_100, n_101, n_102, n_111, n_112, n_113;
  wire n_114, n_115, n_117, n_118, n_119, n_120, n_122, n_123;
  wire n_124, n_125, n_126, n_127, n_128, n_130, n_131, n_132;
  wire n_133, n_135, n_136, n_137, n_138, n_140, n_141, n_142;
  wire n_143, n_145, n_146, n_147, n_148, n_150, n_151, n_152;
  wire n_153, n_155, n_156, n_157, n_158, n_160, n_161, n_162;
  wire n_163, n_164, n_165, n_166, n_167, n_168, n_169, n_170;
  wire n_171;
  xor g15 (n_65, in_0[1], in_2[1]);
  and g16 (n_53, in_0[1], in_2[1]);
  xor g17 (n_73, in_0[2], in_1[2]);
  xor g18 (n_64, n_73, in_2[2]);
  nand g19 (n_74, in_0[2], in_1[2]);
  nand g4 (n_75, in_2[2], in_1[2]);
  nand g5 (n_76, in_0[2], in_2[2]);
  nand g20 (n_52, n_74, n_75, n_76);
  xor g21 (n_77, in_0[3], in_1[3]);
  xor g22 (n_63, n_77, in_2[3]);
  nand g23 (n_78, in_0[3], in_1[3]);
  nand g24 (n_79, in_2[3], in_1[3]);
  nand g25 (n_80, in_0[3], in_2[3]);
  nand g6 (n_51, n_78, n_79, n_80);
  xor g26 (n_66, in_0[4], in_1[4]);
  xor g27 (n_62, n_66, in_2[4]);
  nand g28 (n_67, in_0[4], in_1[4]);
  nand g29 (n_81, in_2[4], in_1[4]);
  nand g30 (n_82, in_0[4], in_2[4]);
  nand g31 (n_50, n_67, n_81, n_82);
  xor g32 (n_83, in_0[5], in_1[5]);
  xor g33 (n_61, n_83, in_2[5]);
  nand g34 (n_84, in_0[5], in_1[5]);
  nand g35 (n_85, in_2[5], in_1[5]);
  nand g36 (n_86, in_0[5], in_2[5]);
  nand g37 (n_49, n_84, n_85, n_86);
  xor g38 (n_87, in_0[6], in_1[6]);
  xor g39 (n_60, n_87, in_2[6]);
  nand g40 (n_88, in_0[6], in_1[6]);
  nand g41 (n_89, in_2[6], in_1[6]);
  nand g42 (n_90, in_0[6], in_2[6]);
  nand g43 (n_48, n_88, n_89, n_90);
  xor g44 (n_91, in_0[7], in_1[7]);
  xor g45 (n_59, n_91, in_2[7]);
  nand g46 (n_92, in_0[7], in_1[7]);
  nand g47 (n_93, in_2[7], in_1[7]);
  nand g48 (n_94, in_0[7], in_2[7]);
  nand g49 (n_47, n_92, n_93, n_94);
  xor g50 (n_95, in_0[8], in_1[8]);
  xor g51 (n_58, n_95, in_2[8]);
  nand g52 (n_96, in_0[8], in_1[8]);
  nand g53 (n_97, in_2[8], in_1[8]);
  nand g54 (n_98, in_0[8], in_2[8]);
  nand g55 (n_46, n_96, n_97, n_98);
  xor g56 (n_99, in_0[9], in_1[9]);
  xor g57 (n_57, n_99, in_2[9]);
  nand g58 (n_100, in_0[9], in_1[9]);
  nand g59 (n_101, in_2[9], in_1[9]);
  nand g60 (n_102, in_0[9], in_2[9]);
  nand g61 (n_45, n_100, n_101, n_102);
  xor g65 (n_56, in_2[10], n_72);
  xor g72 (n_171, in_2[0], in_1[0]);
  nand g73 (n_111, in_2[0], in_1[0]);
  nand g74 (n_112, in_2[0], in_0[0]);
  nand g7 (n_113, in_1[0], in_0[0]);
  nand g8 (n_115, n_111, n_112, n_113);
  nor g9 (n_114, in_1[1], n_65);
  nand g10 (n_117, in_1[1], n_65);
  nor g11 (n_119, n_53, n_64);
  nand g12 (n_122, n_53, n_64);
  nor g13 (n_124, n_52, n_63);
  nand g14 (n_55, n_52, n_63);
  nor g75 (n_127, n_51, n_62);
  nand g76 (n_130, n_51, n_62);
  nor g77 (n_132, n_50, n_61);
  nand g78 (n_135, n_50, n_61);
  nor g79 (n_137, n_49, n_60);
  nand g80 (n_140, n_49, n_60);
  nor g81 (n_142, n_48, n_59);
  nand g82 (n_145, n_48, n_59);
  nor g83 (n_147, n_47, n_58);
  nand g84 (n_150, n_47, n_58);
  nor g85 (n_152, n_46, n_57);
  nand g86 (n_155, n_46, n_57);
  nand g91 (n_120, n_117, n_118);
  nand g94 (n_125, n_122, n_123);
  nand g97 (n_128, n_55, n_126);
  nand g100 (n_133, n_130, n_131);
  nand g103 (n_138, n_135, n_136);
  nand g106 (n_143, n_140, n_141);
  nand g109 (n_148, n_145, n_146);
  nand g112 (n_153, n_150, n_151);
  nand g115 (n_158, n_155, n_156);
  xnor g118 (out_0[1], n_115, n_161);
  xnor g120 (out_0[2], n_120, n_162);
  xnor g122 (out_0[3], n_125, n_163);
  xnor g124 (out_0[4], n_128, n_164);
  xnor g126 (out_0[5], n_133, n_165);
  xnor g128 (out_0[6], n_138, n_166);
  xnor g130 (out_0[7], n_143, n_167);
  xnor g132 (out_0[8], n_148, n_168);
  xnor g134 (out_0[9], n_153, n_169);
  xnor g136 (out_0[10], n_158, n_170);
  xor g137 (out_0[0], in_0[0], n_171);
  xor g138 (n_72, in_0[10], in_1[10]);
  or g139 (n_118, n_114, wc);
  not gc (wc, n_115);
  or g140 (n_161, wc0, n_114);
  not gc0 (wc0, n_117);
  and g141 (n_157, n_45, n_56);
  or g142 (n_160, n_45, n_56);
  or g143 (n_162, wc1, n_119);
  not gc1 (wc1, n_122);
  or g144 (n_163, wc2, n_124);
  not gc2 (wc2, n_55);
  or g145 (n_164, wc3, n_127);
  not gc3 (wc3, n_130);
  or g146 (n_165, wc4, n_132);
  not gc4 (wc4, n_135);
  or g147 (n_166, wc5, n_137);
  not gc5 (wc5, n_140);
  or g148 (n_167, wc6, n_142);
  not gc6 (wc6, n_145);
  or g149 (n_168, wc7, n_147);
  not gc7 (wc7, n_150);
  or g150 (n_169, wc8, n_152);
  not gc8 (wc8, n_155);
  or g151 (n_123, wc9, n_119);
  not gc9 (wc9, n_120);
  or g152 (n_170, wc10, n_157);
  not gc10 (wc10, n_160);
  or g153 (n_126, wc11, n_124);
  not gc11 (wc11, n_125);
  or g154 (n_131, wc12, n_127);
  not gc12 (wc12, n_128);
  or g155 (n_136, wc13, n_132);
  not gc13 (wc13, n_133);
  or g156 (n_141, wc14, n_137);
  not gc14 (wc14, n_138);
  or g157 (n_146, wc15, n_142);
  not gc15 (wc15, n_143);
  or g158 (n_151, wc16, n_147);
  not gc16 (wc16, n_148);
  or g159 (n_156, wc17, n_152);
  not gc17 (wc17, n_153);
endmodule

module csa_tree_add_52_27_group_97_GENERIC(in_0, in_1, in_2, out_0);
  input [10:0] in_0, in_1, in_2;
  output [10:0] out_0;
  wire [10:0] in_0, in_1, in_2;
  wire [10:0] out_0;
  csa_tree_add_52_27_group_97_GENERIC_REAL g1(.in_0 (in_0), .in_1
       (in_1), .in_2 (in_2), .out_0 (out_0));
endmodule

module mult_signed_43_152_GENERIC_REAL(A, B, Z);
// synthesis_equation "assign Z = $signed(A) * $signed(B);"
  input [1:0] A;
  input [9:0] B;
  output [10:0] Z;
  wire [1:0] A;
  wire [9:0] B;
  wire [10:0] Z;
  wire n_25, n_26, n_27, n_28, n_29, n_30, n_31, n_32;
  wire n_33, n_44, n_50, n_54, n_55, n_59, n_60, n_61;
  wire n_62, n_63, n_64, n_65, n_66, n_67, n_68, n_69;
  wire n_70, n_71, n_72, n_73, n_74, n_75, n_76, n_77;
  wire n_78, n_79, n_80, n_81, n_82, n_83, n_84, n_85;
  wire n_88, n_89, n_100, n_103, n_109, n_114, n_119, n_124;
  wire n_129, n_134, n_139, n_144, n_149;
  xor g2 (n_50, A[1], A[0]);
  xor g8 (n_54, A[1], B[0]);
  and g12 (Z[0], B[0], A[0]);
  xor g13 (n_59, A[1], B[1]);
  nand g14 (n_60, n_59, A[0]);
  nand g15 (n_61, n_54, n_55);
  nand g16 (n_44, n_60, n_61);
  xor g17 (n_62, A[1], B[2]);
  nand g18 (n_63, n_62, A[0]);
  nand g19 (n_64, n_59, n_55);
  nand g20 (n_32, n_63, n_64);
  xor g21 (n_65, A[1], B[3]);
  nand g22 (n_66, n_65, A[0]);
  nand g23 (n_67, n_62, n_55);
  nand g24 (n_31, n_66, n_67);
  xor g25 (n_68, A[1], B[4]);
  nand g26 (n_69, n_68, A[0]);
  nand g27 (n_70, n_65, n_55);
  nand g28 (n_30, n_69, n_70);
  xor g29 (n_71, A[1], B[5]);
  nand g30 (n_72, n_71, A[0]);
  nand g31 (n_73, n_68, n_55);
  nand g32 (n_29, n_72, n_73);
  xor g33 (n_74, A[1], B[6]);
  nand g34 (n_75, n_74, A[0]);
  nand g35 (n_76, n_71, n_55);
  nand g36 (n_28, n_75, n_76);
  xor g37 (n_77, A[1], B[7]);
  nand g38 (n_78, n_77, A[0]);
  nand g39 (n_79, n_74, n_55);
  nand g40 (n_27, n_78, n_79);
  xor g41 (n_80, A[1], B[8]);
  nand g42 (n_81, n_80, A[0]);
  nand g43 (n_82, n_77, n_55);
  nand g44 (n_26, n_81, n_82);
  xor g45 (n_83, A[1], B[9]);
  nand g46 (n_84, n_83, A[0]);
  nand g47 (n_85, n_80, n_55);
  nand g48 (n_25, n_84, n_85);
  nand g51 (n_88, n_83, n_55);
  nand g52 (n_89, n_84, n_88);
  nor g65 (n_100, n_33, n_44);
  nand g66 (n_103, n_33, n_44);
  and g135 (n_55, wc, n_50);
  not gc (wc, A[0]);
  and g137 (n_33, A[1], wc0);
  not gc0 (wc0, Z[0]);
  or g147 (n_149, wc1, n_100);
  not gc1 (wc1, n_103);
  not g158 (Z[1], n_149);
  or g159 (n_109, n_103, wc2);
  not gc2 (wc2, n_32);
  xnor g160 (Z[2], n_32, n_103);
  or g162 (n_114, n_109, wc3);
  not gc3 (wc3, n_31);
  xnor g163 (Z[3], n_31, n_109);
  or g165 (n_119, n_114, wc4);
  not gc4 (wc4, n_30);
  xnor g166 (Z[4], n_30, n_114);
  or g168 (n_124, n_119, wc5);
  not gc5 (wc5, n_29);
  xnor g169 (Z[5], n_29, n_119);
  or g171 (n_129, n_124, wc6);
  not gc6 (wc6, n_28);
  xnor g172 (Z[6], n_28, n_124);
  or g174 (n_134, n_129, wc7);
  not gc7 (wc7, n_27);
  xnor g175 (Z[7], n_27, n_129);
  or g177 (n_139, n_134, wc8);
  not gc8 (wc8, n_26);
  xnor g178 (Z[8], n_26, n_134);
  or g180 (n_144, n_139, wc9);
  not gc9 (wc9, n_25);
  xnor g181 (Z[9], n_25, n_139);
  xnor g183 (Z[10], n_89, n_144);
endmodule

module mult_signed_43_152_GENERIC(A, B, Z);
  input [1:0] A;
  input [9:0] B;
  output [10:0] Z;
  wire [1:0] A;
  wire [9:0] B;
  wire [10:0] Z;
  mult_signed_43_152_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module mult_signed_43_GENERIC_REAL(A, B, Z);
// synthesis_equation "assign Z = $signed(A) * $signed(B);"
  input [1:0] A;
  input [9:0] B;
  output [10:0] Z;
  wire [1:0] A;
  wire [9:0] B;
  wire [10:0] Z;
  wire n_25, n_26, n_27, n_28, n_29, n_30, n_31, n_32;
  wire n_33, n_44, n_50, n_54, n_55, n_59, n_60, n_61;
  wire n_62, n_63, n_64, n_65, n_66, n_67, n_68, n_69;
  wire n_70, n_71, n_72, n_73, n_74, n_75, n_76, n_77;
  wire n_78, n_79, n_80, n_81, n_82, n_83, n_84, n_85;
  wire n_88, n_89, n_100, n_103, n_109, n_114, n_119, n_124;
  wire n_129, n_134, n_139, n_144, n_149;
  xor g2 (n_50, A[1], A[0]);
  xor g8 (n_54, A[1], B[0]);
  and g12 (Z[0], B[0], A[0]);
  xor g13 (n_59, A[1], B[1]);
  nand g14 (n_60, n_59, A[0]);
  nand g15 (n_61, n_54, n_55);
  nand g16 (n_44, n_60, n_61);
  xor g17 (n_62, A[1], B[2]);
  nand g18 (n_63, n_62, A[0]);
  nand g19 (n_64, n_59, n_55);
  nand g20 (n_32, n_63, n_64);
  xor g21 (n_65, A[1], B[3]);
  nand g22 (n_66, n_65, A[0]);
  nand g23 (n_67, n_62, n_55);
  nand g24 (n_31, n_66, n_67);
  xor g25 (n_68, A[1], B[4]);
  nand g26 (n_69, n_68, A[0]);
  nand g27 (n_70, n_65, n_55);
  nand g28 (n_30, n_69, n_70);
  xor g29 (n_71, A[1], B[5]);
  nand g30 (n_72, n_71, A[0]);
  nand g31 (n_73, n_68, n_55);
  nand g32 (n_29, n_72, n_73);
  xor g33 (n_74, A[1], B[6]);
  nand g34 (n_75, n_74, A[0]);
  nand g35 (n_76, n_71, n_55);
  nand g36 (n_28, n_75, n_76);
  xor g37 (n_77, A[1], B[7]);
  nand g38 (n_78, n_77, A[0]);
  nand g39 (n_79, n_74, n_55);
  nand g40 (n_27, n_78, n_79);
  xor g41 (n_80, A[1], B[8]);
  nand g42 (n_81, n_80, A[0]);
  nand g43 (n_82, n_77, n_55);
  nand g44 (n_26, n_81, n_82);
  xor g45 (n_83, A[1], B[9]);
  nand g46 (n_84, n_83, A[0]);
  nand g47 (n_85, n_80, n_55);
  nand g48 (n_25, n_84, n_85);
  nand g51 (n_88, n_83, n_55);
  nand g52 (n_89, n_84, n_88);
  nor g65 (n_100, n_33, n_44);
  nand g66 (n_103, n_33, n_44);
  and g135 (n_55, wc, n_50);
  not gc (wc, A[0]);
  and g137 (n_33, A[1], wc0);
  not gc0 (wc0, Z[0]);
  or g147 (n_149, wc1, n_100);
  not gc1 (wc1, n_103);
  not g158 (Z[1], n_149);
  or g159 (n_109, n_103, wc2);
  not gc2 (wc2, n_32);
  xnor g160 (Z[2], n_32, n_103);
  or g162 (n_114, n_109, wc3);
  not gc3 (wc3, n_31);
  xnor g163 (Z[3], n_31, n_109);
  or g165 (n_119, n_114, wc4);
  not gc4 (wc4, n_30);
  xnor g166 (Z[4], n_30, n_114);
  or g168 (n_124, n_119, wc5);
  not gc5 (wc5, n_29);
  xnor g169 (Z[5], n_29, n_119);
  or g171 (n_129, n_124, wc6);
  not gc6 (wc6, n_28);
  xnor g172 (Z[6], n_28, n_124);
  or g174 (n_134, n_129, wc7);
  not gc7 (wc7, n_27);
  xnor g175 (Z[7], n_27, n_129);
  or g177 (n_139, n_134, wc8);
  not gc8 (wc8, n_26);
  xnor g178 (Z[8], n_26, n_134);
  or g180 (n_144, n_139, wc9);
  not gc9 (wc9, n_25);
  xnor g181 (Z[9], n_25, n_139);
  xnor g183 (Z[10], n_89, n_144);
endmodule

module mult_signed_43_GENERIC(A, B, Z);
  input [1:0] A;
  input [9:0] B;
  output [10:0] Z;
  wire [1:0] A;
  wire [9:0] B;
  wire [10:0] Z;
  mult_signed_43_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module mult_signed_43_153_GENERIC_REAL(A, B, Z);
// synthesis_equation "assign Z = $signed(A) * $signed(B);"
  input [1:0] A;
  input [9:0] B;
  output [10:0] Z;
  wire [1:0] A;
  wire [9:0] B;
  wire [10:0] Z;
  wire n_25, n_26, n_27, n_28, n_29, n_30, n_31, n_32;
  wire n_33, n_44, n_50, n_54, n_55, n_59, n_60, n_61;
  wire n_62, n_63, n_64, n_65, n_66, n_67, n_68, n_69;
  wire n_70, n_71, n_72, n_73, n_74, n_75, n_76, n_77;
  wire n_78, n_79, n_80, n_81, n_82, n_83, n_84, n_85;
  wire n_88, n_89, n_100, n_103, n_109, n_114, n_119, n_124;
  wire n_129, n_134, n_139, n_144, n_149;
  xor g2 (n_50, A[1], A[0]);
  xor g8 (n_54, A[1], B[0]);
  and g12 (Z[0], B[0], A[0]);
  xor g13 (n_59, A[1], B[1]);
  nand g14 (n_60, n_59, A[0]);
  nand g15 (n_61, n_54, n_55);
  nand g16 (n_44, n_60, n_61);
  xor g17 (n_62, A[1], B[2]);
  nand g18 (n_63, n_62, A[0]);
  nand g19 (n_64, n_59, n_55);
  nand g20 (n_32, n_63, n_64);
  xor g21 (n_65, A[1], B[3]);
  nand g22 (n_66, n_65, A[0]);
  nand g23 (n_67, n_62, n_55);
  nand g24 (n_31, n_66, n_67);
  xor g25 (n_68, A[1], B[4]);
  nand g26 (n_69, n_68, A[0]);
  nand g27 (n_70, n_65, n_55);
  nand g28 (n_30, n_69, n_70);
  xor g29 (n_71, A[1], B[5]);
  nand g30 (n_72, n_71, A[0]);
  nand g31 (n_73, n_68, n_55);
  nand g32 (n_29, n_72, n_73);
  xor g33 (n_74, A[1], B[6]);
  nand g34 (n_75, n_74, A[0]);
  nand g35 (n_76, n_71, n_55);
  nand g36 (n_28, n_75, n_76);
  xor g37 (n_77, A[1], B[7]);
  nand g38 (n_78, n_77, A[0]);
  nand g39 (n_79, n_74, n_55);
  nand g40 (n_27, n_78, n_79);
  xor g41 (n_80, A[1], B[8]);
  nand g42 (n_81, n_80, A[0]);
  nand g43 (n_82, n_77, n_55);
  nand g44 (n_26, n_81, n_82);
  xor g45 (n_83, A[1], B[9]);
  nand g46 (n_84, n_83, A[0]);
  nand g47 (n_85, n_80, n_55);
  nand g48 (n_25, n_84, n_85);
  nand g51 (n_88, n_83, n_55);
  nand g52 (n_89, n_84, n_88);
  nor g65 (n_100, n_33, n_44);
  nand g66 (n_103, n_33, n_44);
  and g135 (n_55, wc, n_50);
  not gc (wc, A[0]);
  and g137 (n_33, A[1], wc0);
  not gc0 (wc0, Z[0]);
  or g147 (n_149, wc1, n_100);
  not gc1 (wc1, n_103);
  not g158 (Z[1], n_149);
  or g159 (n_109, n_103, wc2);
  not gc2 (wc2, n_32);
  xnor g160 (Z[2], n_32, n_103);
  or g162 (n_114, n_109, wc3);
  not gc3 (wc3, n_31);
  xnor g163 (Z[3], n_31, n_109);
  or g165 (n_119, n_114, wc4);
  not gc4 (wc4, n_30);
  xnor g166 (Z[4], n_30, n_114);
  or g168 (n_124, n_119, wc5);
  not gc5 (wc5, n_29);
  xnor g169 (Z[5], n_29, n_119);
  or g171 (n_129, n_124, wc6);
  not gc6 (wc6, n_28);
  xnor g172 (Z[6], n_28, n_124);
  or g174 (n_134, n_129, wc7);
  not gc7 (wc7, n_27);
  xnor g175 (Z[7], n_27, n_129);
  or g177 (n_139, n_134, wc8);
  not gc8 (wc8, n_26);
  xnor g178 (Z[8], n_26, n_134);
  or g180 (n_144, n_139, wc9);
  not gc9 (wc9, n_25);
  xnor g181 (Z[9], n_25, n_139);
  xnor g183 (Z[10], n_89, n_144);
endmodule

module mult_signed_43_153_GENERIC(A, B, Z);
  input [1:0] A;
  input [9:0] B;
  output [10:0] Z;
  wire [1:0] A;
  wire [9:0] B;
  wire [10:0] Z;
  mult_signed_43_153_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

