module csa_tree_add_100_25_group_194_GENERIC_REAL(in_0, in_1, in_2,
     out_0);
// synthesis_equation "assign out_0 = ( $signed(in_2) + ( $signed(in_0) * $signed(in_1) )  )  ;"
  input [8:0] in_0;
  input [1:0] in_1;
  input [15:0] in_2;
  output [15:0] out_0;
  wire [8:0] in_0;
  wire [1:0] in_1;
  wire [15:0] in_2;
  wire [15:0] out_0;
  wire n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57;
  wire n_58, n_59, n_65, n_66, n_67, n_68, n_69, n_70;
  wire n_71, n_72, n_73, n_74, n_76, n_78, n_79, n_80;
  wire n_81, n_82, n_83, n_84, n_85, n_86, n_87, n_88;
  wire n_89, n_90, n_92, n_93, n_95, n_105, n_106, n_107;
  wire n_108, n_109, n_110, n_111, n_112, n_113, n_114, n_115;
  wire n_116, n_117, n_118, n_119, n_120, n_121, n_122, n_123;
  wire n_124, n_125, n_126, n_127, n_128, n_129, n_130, n_131;
  wire n_132, n_133, n_134, n_135, n_136, n_137, n_141, n_143;
  wire n_146, n_147, n_148, n_149, n_151, n_152, n_153, n_154;
  wire n_156, n_157, n_158, n_159, n_161, n_162, n_163, n_165;
  wire n_166, n_167, n_168, n_170, n_171, n_172, n_173, n_175;
  wire n_176, n_177, n_178, n_180, n_181, n_182, n_183, n_185;
  wire n_186, n_187, n_188, n_190, n_191, n_192, n_193, n_195;
  wire n_196, n_197, n_198, n_200, n_201, n_202, n_203, n_205;
  wire n_206, n_207, n_208, n_210, n_211, n_212, n_213, n_215;
  wire n_216, n_217, n_218, n_219, n_220, n_221, n_222, n_223;
  wire n_224, n_225, n_226, n_227, n_228, n_229, n_230;
  and g2 (n_59, in_0[0], in_1[0]);
  and g3 (n_58, in_0[1], in_1[0]);
  and g4 (n_79, in_0[2], in_1[0]);
  and g5 (n_81, in_0[3], in_1[0]);
  and g6 (n_83, in_0[4], in_1[0]);
  and g7 (n_85, in_0[5], in_1[0]);
  and g8 (n_87, in_0[6], in_1[0]);
  and g9 (n_89, in_0[7], in_1[0]);
  nand g10 (n_92, in_0[8], in_1[0]);
  nand g11 (n_78, in_0[0], in_1[1]);
  nand g12 (n_80, in_0[1], in_1[1]);
  nand g13 (n_82, in_0[2], in_1[1]);
  nand g14 (n_84, in_0[3], in_1[1]);
  nand g15 (n_86, in_0[4], in_1[1]);
  nand g16 (n_88, in_0[5], in_1[1]);
  nand g17 (n_90, in_0[6], in_1[1]);
  nand g18 (n_93, in_0[7], in_1[1]);
  and g19 (n_95, in_0[8], in_1[1]);
  nand g39 (n_105, in_2[1], n_78);
  xor g41 (n_106, in_2[2], n_79);
  xor g42 (n_73, n_106, n_80);
  nand g43 (n_107, in_2[2], n_79);
  nand g44 (n_108, n_80, n_79);
  nand g45 (n_109, in_2[2], n_80);
  nand g46 (n_56, n_107, n_108, n_109);
  xor g47 (n_110, in_2[3], n_81);
  xor g48 (n_72, n_110, n_82);
  nand g49 (n_111, in_2[3], n_81);
  nand g50 (n_112, n_82, n_81);
  nand g51 (n_113, in_2[3], n_82);
  nand g52 (n_55, n_111, n_112, n_113);
  xor g53 (n_114, in_2[4], n_83);
  xor g54 (n_71, n_114, n_84);
  nand g55 (n_115, in_2[4], n_83);
  nand g56 (n_116, n_84, n_83);
  nand g57 (n_117, in_2[4], n_84);
  nand g58 (n_54, n_115, n_116, n_117);
  xor g59 (n_118, in_2[5], n_85);
  xor g60 (n_70, n_118, n_86);
  nand g61 (n_119, in_2[5], n_85);
  nand g62 (n_120, n_86, n_85);
  nand g63 (n_121, in_2[5], n_86);
  nand g64 (n_53, n_119, n_120, n_121);
  xor g65 (n_122, in_2[6], n_87);
  xor g66 (n_69, n_122, n_88);
  nand g67 (n_123, in_2[6], n_87);
  nand g68 (n_124, n_88, n_87);
  nand g69 (n_125, in_2[6], n_88);
  nand g70 (n_52, n_123, n_124, n_125);
  xor g71 (n_126, in_2[7], n_89);
  xor g72 (n_68, n_126, n_90);
  nand g73 (n_127, in_2[7], n_89);
  nand g74 (n_128, n_90, n_89);
  nand g75 (n_129, in_2[7], n_90);
  nand g76 (n_51, n_127, n_128, n_129);
  xor g79 (n_130, n_92, n_93);
  nand g81 (n_131, n_92, n_93);
  nand g84 (n_50, n_131, n_132, n_133);
  xor g85 (n_134, in_2[9], n_95);
  xor g86 (n_66, n_134, in_2[8]);
  nand g87 (n_135, in_2[9], n_95);
  nand g88 (n_136, in_2[8], n_95);
  nand g89 (n_137, in_2[9], in_2[8]);
  nand g90 (n_65, n_135, n_136, n_137);
  nand g105 (n_141, n_59, in_2[0]);
  nor g108 (n_143, n_58, n_74);
  nand g109 (n_146, n_58, n_74);
  nor g110 (n_148, n_57, n_73);
  nand g111 (n_151, n_57, n_73);
  nor g112 (n_153, n_56, n_72);
  nand g113 (n_156, n_56, n_72);
  nor g114 (n_158, n_55, n_71);
  nand g115 (n_161, n_55, n_71);
  nor g116 (n_162, n_54, n_70);
  nand g117 (n_165, n_54, n_70);
  nor g118 (n_167, n_53, n_69);
  nand g20 (n_170, n_53, n_69);
  nor g21 (n_172, n_52, n_68);
  nand g22 (n_175, n_52, n_68);
  nor g23 (n_177, n_51, n_67);
  nand g24 (n_180, n_51, n_67);
  nor g25 (n_182, n_50, n_66);
  nand g26 (n_185, n_50, n_66);
  nand g125 (n_149, n_146, n_147);
  nand g128 (n_154, n_151, n_152);
  nand g131 (n_159, n_156, n_157);
  nand g134 (n_163, n_161, n_76);
  nand g137 (n_168, n_165, n_166);
  nand g140 (n_173, n_170, n_171);
  nand g143 (n_178, n_175, n_176);
  nand g146 (n_183, n_180, n_181);
  nand g149 (n_188, n_185, n_186);
  nand g152 (n_193, n_190, n_191);
  nand g155 (n_198, n_195, n_196);
  nand g158 (n_203, n_200, n_201);
  nand g161 (n_208, n_205, n_206);
  nand g164 (n_213, n_210, n_211);
  xnor g169 (out_0[2], n_149, n_217);
  xnor g171 (out_0[3], n_154, n_218);
  xnor g173 (out_0[4], n_159, n_219);
  xnor g175 (out_0[5], n_163, n_220);
  xnor g177 (out_0[6], n_168, n_221);
  xnor g179 (out_0[7], n_173, n_222);
  xnor g181 (out_0[8], n_178, n_223);
  xnor g183 (out_0[9], n_183, n_224);
  xnor g185 (out_0[10], n_188, n_225);
  xnor g187 (out_0[11], n_193, n_226);
  xnor g189 (out_0[12], n_198, n_227);
  xnor g191 (out_0[13], n_203, n_228);
  xnor g193 (out_0[14], n_208, n_229);
  xnor g195 (out_0[15], n_213, n_230);
  xor g196 (out_0[0], in_2[0], n_59);
  xnor g204 (n_74, n_78, in_2[1]);
  or g206 (n_132, in_2[8], wc);
  not gc (wc, n_93);
  or g207 (n_133, in_2[8], wc0);
  not gc0 (wc0, n_92);
  and g208 (n_192, wc1, in_2[11]);
  not gc1 (wc1, in_2[10]);
  or g209 (n_195, wc2, in_2[11]);
  not gc2 (wc2, in_2[10]);
  and g210 (n_197, wc3, in_2[12]);
  not gc3 (wc3, in_2[11]);
  or g211 (n_200, wc4, in_2[12]);
  not gc4 (wc4, in_2[11]);
  and g212 (n_202, wc5, in_2[13]);
  not gc5 (wc5, in_2[12]);
  or g213 (n_205, wc6, in_2[13]);
  not gc6 (wc6, in_2[12]);
  and g214 (n_207, wc7, in_2[14]);
  not gc7 (wc7, in_2[13]);
  or g215 (n_210, wc8, in_2[14]);
  not gc8 (wc8, in_2[13]);
  or g216 (n_57, in_2[1], wc9, n_78);
  not gc9 (wc9, n_105);
  xnor g217 (n_67, n_130, in_2[8]);
  and g219 (n_212, in_2[14], wc10);
  not gc10 (wc10, in_2[15]);
  or g220 (n_215, in_2[14], wc11);
  not gc11 (wc11, in_2[15]);
  and g221 (n_187, in_2[10], wc12);
  not gc12 (wc12, n_65);
  or g222 (n_190, in_2[10], wc13);
  not gc13 (wc13, n_65);
  or g223 (n_226, wc14, n_192);
  not gc14 (wc14, n_195);
  or g224 (n_227, wc15, n_197);
  not gc15 (wc15, n_200);
  or g225 (n_228, wc16, n_202);
  not gc16 (wc16, n_205);
  or g226 (n_229, wc17, n_207);
  not gc17 (wc17, n_210);
  or g227 (n_147, n_141, n_143);
  or g228 (n_216, wc18, n_143);
  not gc18 (wc18, n_146);
  or g229 (n_230, wc19, n_212);
  not gc19 (wc19, n_215);
  xor g230 (out_0[1], n_141, n_216);
  or g231 (n_217, wc20, n_148);
  not gc20 (wc20, n_151);
  or g232 (n_218, wc21, n_153);
  not gc21 (wc21, n_156);
  or g233 (n_219, wc22, n_158);
  not gc22 (wc22, n_161);
  or g234 (n_220, wc23, n_162);
  not gc23 (wc23, n_165);
  or g235 (n_221, wc24, n_167);
  not gc24 (wc24, n_170);
  or g236 (n_222, wc25, n_172);
  not gc25 (wc25, n_175);
  or g237 (n_223, wc26, n_177);
  not gc26 (wc26, n_180);
  or g238 (n_224, wc27, n_182);
  not gc27 (wc27, n_185);
  or g239 (n_225, wc28, n_187);
  not gc28 (wc28, n_190);
  or g240 (n_152, wc29, n_148);
  not gc29 (wc29, n_149);
  or g241 (n_157, wc30, n_153);
  not gc30 (wc30, n_154);
  or g242 (n_76, wc31, n_158);
  not gc31 (wc31, n_159);
  or g243 (n_166, wc32, n_162);
  not gc32 (wc32, n_163);
  or g244 (n_171, wc33, n_167);
  not gc33 (wc33, n_168);
  or g245 (n_176, wc34, n_172);
  not gc34 (wc34, n_173);
  or g246 (n_181, wc35, n_177);
  not gc35 (wc35, n_178);
  or g247 (n_186, wc36, n_182);
  not gc36 (wc36, n_183);
  or g248 (n_191, n_187, wc37);
  not gc37 (wc37, n_188);
  or g249 (n_196, n_192, wc38);
  not gc38 (wc38, n_193);
  or g250 (n_201, n_197, wc39);
  not gc39 (wc39, n_198);
  or g251 (n_206, n_202, wc40);
  not gc40 (wc40, n_203);
  or g252 (n_211, n_207, wc41);
  not gc41 (wc41, n_208);
endmodule

module csa_tree_add_100_25_group_194_GENERIC(in_0, in_1, in_2, out_0);
  input [8:0] in_0;
  input [1:0] in_1;
  input [15:0] in_2;
  output [15:0] out_0;
  wire [8:0] in_0;
  wire [1:0] in_1;
  wire [15:0] in_2;
  wire [15:0] out_0;
  csa_tree_add_100_25_group_194_GENERIC_REAL g1(.in_0 (in_0), .in_1
       (in_1), .in_2 (in_2), .out_0 (out_0));
endmodule

