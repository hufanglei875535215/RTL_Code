module csa_tree_add_64_12_group_14_GENERIC_REAL(in_0, in_1, in_2,
     out_0);
// synthesis_equation "assign out_0 = ( $signed(in_2) + ( $signed(in_0) * $signed(in_1) )  )  ;"
  input [1:0] in_0;
  input [8:0] in_1, in_2;
  output [8:0] out_0;
  wire [1:0] in_0;
  wire [8:0] in_1, in_2;
  wire [8:0] out_0;
  wire n_30, n_31, n_32, n_33, n_34, n_35, n_36, n_37;
  wire n_38, n_39, n_40, n_41, n_42, n_43, n_44, n_45;
  wire n_46, n_48, n_52, n_56, n_57, n_61, n_62, n_63;
  wire n_64, n_65, n_66, n_67, n_68, n_69, n_70, n_71;
  wire n_72, n_73, n_74, n_75, n_76, n_77, n_78, n_79;
  wire n_80, n_81, n_82, n_83, n_89, n_90, n_91, n_92;
  wire n_93, n_94, n_95, n_98, n_107, n_109, n_112, n_113;
  wire n_114, n_115, n_117, n_118, n_119, n_120, n_122, n_123;
  wire n_124, n_125, n_127, n_128, n_129, n_130, n_132, n_133;
  wire n_134, n_135, n_137, n_138, n_139, n_140, n_142, n_143;
  wire n_144, n_145, n_147, n_148, n_149, n_150, n_151, n_152;
  wire n_153, n_154, n_155;
  xor g3 (n_52, in_0[1], in_0[0]);
  xor g9 (n_56, in_0[1], in_1[0]);
  and g13 (n_38, in_1[0], in_0[0]);
  xor g14 (n_61, in_0[1], in_1[1]);
  nand g15 (n_62, n_61, in_0[0]);
  nand g16 (n_63, n_56, n_57);
  nand g17 (n_37, n_62, n_63);
  xor g18 (n_64, in_0[1], in_1[2]);
  nand g19 (n_65, n_64, in_0[0]);
  nand g20 (n_66, n_61, n_57);
  nand g21 (n_36, n_65, n_66);
  xor g22 (n_67, in_0[1], in_1[3]);
  nand g23 (n_68, n_67, in_0[0]);
  nand g24 (n_69, n_64, n_57);
  nand g25 (n_91, n_68, n_69);
  xor g26 (n_70, in_0[1], in_1[4]);
  nand g27 (n_71, n_70, in_0[0]);
  nand g28 (n_72, n_67, n_57);
  nand g29 (n_92, n_71, n_72);
  xor g30 (n_73, in_0[1], in_1[5]);
  nand g31 (n_74, n_73, in_0[0]);
  nand g32 (n_75, n_70, n_57);
  nand g33 (n_93, n_74, n_75);
  xor g34 (n_76, in_0[1], in_1[6]);
  nand g35 (n_77, n_76, in_0[0]);
  nand g36 (n_78, n_73, n_57);
  nand g37 (n_94, n_77, n_78);
  xor g38 (n_79, in_0[1], in_1[7]);
  nand g39 (n_80, n_79, in_0[0]);
  nand g40 (n_81, n_76, n_57);
  nand g41 (n_95, n_80, n_81);
  xor g42 (n_82, in_0[1], in_1[8]);
  nand g43 (n_83, n_82, in_0[0]);
  nand g44 (n_48, n_79, n_57);
  nand g45 (n_98, n_83, n_48);
  xor g58 (n_46, in_2[1], n_89);
  and g59 (n_90, in_2[1], n_89);
  xor g60 (n_45, in_2[2], n_90);
  and g61 (n_35, in_2[2], n_90);
  xor g62 (n_44, in_2[3], n_91);
  and g63 (n_34, in_2[3], n_91);
  xor g64 (n_43, in_2[4], n_92);
  and g65 (n_33, in_2[4], n_92);
  xor g66 (n_42, in_2[5], n_93);
  and g67 (n_32, in_2[5], n_93);
  xor g68 (n_41, in_2[6], n_94);
  and g69 (n_31, in_2[6], n_94);
  xor g70 (n_40, in_2[7], n_95);
  and g71 (n_30, in_2[7], n_95);
  xor g73 (n_39, in_2[8], n_98);
  nand g82 (n_107, n_38, in_2[0]);
  nor g85 (n_109, n_37, n_46);
  nand g86 (n_112, n_37, n_46);
  nor g87 (n_114, n_36, n_45);
  nand g88 (n_117, n_36, n_45);
  nor g89 (n_119, n_35, n_44);
  nand g90 (n_122, n_35, n_44);
  nor g91 (n_124, n_34, n_43);
  nand g92 (n_127, n_34, n_43);
  nor g93 (n_129, n_33, n_42);
  nand g94 (n_132, n_33, n_42);
  nor g95 (n_134, n_32, n_41);
  nand g96 (n_137, n_32, n_41);
  nor g97 (n_139, n_31, n_40);
  nand g98 (n_142, n_31, n_40);
  nand g103 (n_115, n_112, n_113);
  nand g106 (n_120, n_117, n_118);
  nand g109 (n_125, n_122, n_123);
  nand g112 (n_130, n_127, n_128);
  nand g115 (n_135, n_132, n_133);
  nand g118 (n_140, n_137, n_138);
  nand g121 (n_145, n_142, n_143);
  xnor g52 (out_0[2], n_115, n_149);
  xnor g54 (out_0[3], n_120, n_150);
  xnor g56 (out_0[4], n_125, n_151);
  xnor g124 (out_0[5], n_130, n_152);
  xnor g126 (out_0[6], n_135, n_153);
  xnor g128 (out_0[7], n_140, n_154);
  xnor g130 (out_0[8], n_145, n_155);
  xor g131 (out_0[0], in_2[0], n_38);
  and g133 (n_57, wc, n_52);
  not gc (wc, in_0[0]);
  and g135 (n_89, in_0[1], wc0);
  not gc0 (wc0, n_38);
  and g137 (n_144, n_30, n_39);
  or g138 (n_147, n_30, n_39);
  or g139 (n_113, n_107, n_109);
  or g140 (n_148, wc1, n_109);
  not gc1 (wc1, n_112);
  xor g141 (out_0[1], n_107, n_148);
  or g142 (n_149, wc2, n_114);
  not gc2 (wc2, n_117);
  or g143 (n_150, wc3, n_119);
  not gc3 (wc3, n_122);
  or g144 (n_151, wc4, n_124);
  not gc4 (wc4, n_127);
  or g145 (n_152, wc5, n_129);
  not gc5 (wc5, n_132);
  or g146 (n_153, wc6, n_134);
  not gc6 (wc6, n_137);
  or g147 (n_154, wc7, n_139);
  not gc7 (wc7, n_142);
  or g148 (n_118, wc8, n_114);
  not gc8 (wc8, n_115);
  or g149 (n_155, wc9, n_144);
  not gc9 (wc9, n_147);
  or g150 (n_123, wc10, n_119);
  not gc10 (wc10, n_120);
  or g151 (n_128, wc11, n_124);
  not gc11 (wc11, n_125);
  or g152 (n_133, wc12, n_129);
  not gc12 (wc12, n_130);
  or g153 (n_138, wc13, n_134);
  not gc13 (wc13, n_135);
  or g154 (n_143, wc14, n_139);
  not gc14 (wc14, n_140);
endmodule

module csa_tree_add_64_12_group_14_GENERIC(in_0, in_1, in_2, out_0);
  input [1:0] in_0;
  input [8:0] in_1, in_2;
  output [8:0] out_0;
  wire [1:0] in_0;
  wire [8:0] in_1, in_2;
  wire [8:0] out_0;
  csa_tree_add_64_12_group_14_GENERIC_REAL g1(.in_0 (in_0), .in_1
       (in_1), .in_2 (in_2), .out_0 (out_0));
endmodule

module lt_signed_GENERIC_REAL(A, B, Z);
// synthesis_equation lt_signed
  input [8:0] A;
  input B;
  output Z;
  wire [8:0] A;
  wire B;
  wire Z;
  wire n_32, n_33, n_34, n_35, n_36, n_38, n_39, n_40;
  wire n_43, n_44, n_46, n_47, n_48, n_49, n_50, n_51;
  wire n_53, n_54, n_55, n_57, n_58, n_61, n_62, n_63;
  wire n_64, n_67, n_69, n_71, n_72, n_74, n_82, n_84;
  wire n_85, n_86, n_87, n_89, n_90;
  not g11 (Z, n_39);
  nand g34 (n_58, n_46, n_47);
  nor g35 (n_51, n_48, n_49);
  nor g38 (n_61, n_32, n_49);
  nor g39 (n_36, n_33, n_34);
  nor g42 (n_67, n_38, n_34);
  nor g43 (n_55, n_53, n_40);
  nor g46 (n_69, n_57, n_40);
  nand g50 (n_63, n_61, n_58);
  nand g51 (n_74, n_62, n_63);
  nand g61 (n_82, n_67, n_69);
  nand g72 (n_87, n_84, n_85);
  nand g75 (n_39, n_89, n_90);
  or g98 (n_89, wc, A[8]);
  not gc (wc, B);
  or g99 (n_33, B, wc0);
  not gc0 (wc0, A[4]);
  and g100 (n_34, B, wc1);
  not gc1 (wc1, A[5]);
  or g101 (n_35, B, wc2);
  not gc2 (wc2, A[5]);
  and g102 (n_57, B, wc3);
  not gc3 (wc3, A[6]);
  and g103 (n_40, B, wc4);
  not gc4 (wc4, A[7]);
  or g104 (n_53, B, wc5);
  not gc5 (wc5, A[6]);
  or g105 (n_54, B, wc6);
  not gc6 (wc6, A[7]);
  or g106 (n_48, B, wc7);
  not gc7 (wc7, A[2]);
  and g107 (n_49, B, wc8);
  not gc8 (wc8, A[3]);
  or g108 (n_50, B, wc9);
  not gc9 (wc9, A[3]);
  and g109 (n_32, B, wc10);
  not gc10 (wc10, A[2]);
  or g110 (n_46, B, wc11);
  not gc11 (wc11, A[1]);
  or g111 (n_44, wc12, A[0]);
  not gc12 (wc12, B);
  and g112 (n_43, B, wc13);
  not gc13 (wc13, A[1]);
  and g113 (n_38, B, wc14);
  not gc14 (wc14, A[4]);
  and g114 (n_86, wc15, A[8]);
  not gc15 (wc15, B);
  and g115 (n_64, n_35, wc16);
  not gc16 (wc16, n_36);
  and g116 (n_71, n_54, wc17);
  not gc17 (wc17, n_55);
  and g117 (n_62, n_50, wc18);
  not gc18 (wc18, n_51);
  or g118 (n_47, n_43, wc19);
  not gc19 (wc19, n_44);
  and g119 (n_72, wc20, n_69);
  not gc20 (wc20, n_64);
  and g120 (n_84, wc21, n_71);
  not gc21 (wc21, n_72);
  or g121 (n_85, n_82, wc22);
  not gc22 (wc22, n_74);
  or g122 (n_90, n_86, wc23);
  not gc23 (wc23, n_87);
endmodule

module lt_signed_GENERIC(A, B, Z);
  input [8:0] A;
  input B;
  output Z;
  wire [8:0] A;
  wire B;
  wire Z;
  lt_signed_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

