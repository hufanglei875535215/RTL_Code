module csa_tree_add_133_23_group_102_GENERIC_REAL(in_0, in_1, in_2,
     out_0);
// synthesis_equation "assign out_0 = ( ( $signed(in_1) + $signed(in_2) )  + $signed(in_0) )  ;"
  input [8:0] in_0, in_1, in_2;
  output [8:0] out_0;
  wire [8:0] in_0, in_1, in_2;
  wire [8:0] out_0;
  wire n_37, n_38, n_39, n_40, n_41, n_42, n_43, n_44;
  wire n_45, n_46, n_47, n_48, n_49, n_50, n_51, n_52;
  wire n_53, n_54, n_55, n_60, n_61, n_62, n_63, n_64;
  wire n_65, n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  wire n_73, n_74, n_75, n_76, n_77, n_78, n_79, n_80;
  wire n_81, n_82, n_91, n_92, n_93, n_94, n_95, n_97;
  wire n_98, n_99, n_100, n_102, n_103, n_105, n_106, n_107;
  wire n_108, n_110, n_111, n_112, n_113, n_115, n_116, n_117;
  wire n_118, n_120, n_121, n_122, n_123, n_125, n_126, n_127;
  wire n_128, n_130, n_131, n_132, n_133, n_134, n_135, n_136;
  wire n_137, n_138, n_139;
  xor g13 (n_53, in_0[1], in_2[1]);
  and g14 (n_43, in_0[1], in_2[1]);
  xor g15 (n_61, in_0[2], in_1[2]);
  xor g16 (n_52, n_61, in_2[2]);
  nand g17 (n_62, in_0[2], in_1[2]);
  nand g4 (n_63, in_2[2], in_1[2]);
  nand g5 (n_64, in_0[2], in_2[2]);
  nand g18 (n_42, n_62, n_63, n_64);
  xor g19 (n_65, in_0[3], in_1[3]);
  xor g20 (n_51, n_65, in_2[3]);
  nand g21 (n_66, in_0[3], in_1[3]);
  nand g22 (n_54, in_2[3], in_1[3]);
  nand g23 (n_55, in_0[3], in_2[3]);
  nand g6 (n_41, n_66, n_54, n_55);
  xor g24 (n_67, in_0[4], in_1[4]);
  xor g25 (n_50, n_67, in_2[4]);
  nand g26 (n_68, in_0[4], in_1[4]);
  nand g27 (n_69, in_2[4], in_1[4]);
  nand g28 (n_70, in_0[4], in_2[4]);
  nand g29 (n_40, n_68, n_69, n_70);
  xor g30 (n_71, in_0[5], in_1[5]);
  xor g31 (n_49, n_71, in_2[5]);
  nand g32 (n_72, in_0[5], in_1[5]);
  nand g33 (n_73, in_2[5], in_1[5]);
  nand g34 (n_74, in_0[5], in_2[5]);
  nand g35 (n_39, n_72, n_73, n_74);
  xor g36 (n_75, in_0[6], in_1[6]);
  xor g37 (n_48, n_75, in_2[6]);
  nand g38 (n_76, in_0[6], in_1[6]);
  nand g39 (n_77, in_2[6], in_1[6]);
  nand g40 (n_78, in_0[6], in_2[6]);
  nand g41 (n_38, n_76, n_77, n_78);
  xor g42 (n_79, in_0[7], in_1[7]);
  xor g43 (n_47, n_79, in_2[7]);
  nand g44 (n_80, in_0[7], in_1[7]);
  nand g45 (n_81, in_2[7], in_1[7]);
  nand g46 (n_82, in_0[7], in_2[7]);
  nand g47 (n_37, n_80, n_81, n_82);
  xor g51 (n_46, in_2[8], n_60);
  xor g58 (n_139, in_2[0], in_1[0]);
  nand g59 (n_91, in_2[0], in_1[0]);
  nand g60 (n_92, in_2[0], in_0[0]);
  nand g7 (n_93, in_1[0], in_0[0]);
  nand g8 (n_95, n_91, n_92, n_93);
  nor g9 (n_94, in_1[1], n_53);
  nand g10 (n_97, in_1[1], n_53);
  nor g11 (n_99, n_43, n_52);
  nand g12 (n_44, n_43, n_52);
  nor g61 (n_102, n_42, n_51);
  nand g62 (n_105, n_42, n_51);
  nor g63 (n_107, n_41, n_50);
  nand g64 (n_110, n_41, n_50);
  nor g65 (n_112, n_40, n_49);
  nand g66 (n_115, n_40, n_49);
  nor g67 (n_117, n_39, n_48);
  nand g68 (n_120, n_39, n_48);
  nor g69 (n_122, n_38, n_47);
  nand g70 (n_125, n_38, n_47);
  nand g75 (n_100, n_97, n_98);
  nand g78 (n_103, n_44, n_45);
  nand g81 (n_108, n_105, n_106);
  nand g84 (n_113, n_110, n_111);
  nand g87 (n_118, n_115, n_116);
  nand g90 (n_123, n_120, n_121);
  nand g93 (n_128, n_125, n_126);
  xnor g96 (out_0[1], n_95, n_131);
  xnor g98 (out_0[2], n_100, n_132);
  xnor g100 (out_0[3], n_103, n_133);
  xnor g102 (out_0[4], n_108, n_134);
  xnor g104 (out_0[5], n_113, n_135);
  xnor g106 (out_0[6], n_118, n_136);
  xnor g108 (out_0[7], n_123, n_137);
  xnor g110 (out_0[8], n_128, n_138);
  xor g111 (out_0[0], in_0[0], n_139);
  xor g112 (n_60, in_0[8], in_1[8]);
  or g113 (n_98, n_94, wc);
  not gc (wc, n_95);
  or g114 (n_131, wc0, n_94);
  not gc0 (wc0, n_97);
  and g115 (n_127, n_37, n_46);
  or g116 (n_130, n_37, n_46);
  or g117 (n_132, wc1, n_99);
  not gc1 (wc1, n_44);
  or g118 (n_133, wc2, n_102);
  not gc2 (wc2, n_105);
  or g119 (n_134, wc3, n_107);
  not gc3 (wc3, n_110);
  or g120 (n_135, wc4, n_112);
  not gc4 (wc4, n_115);
  or g121 (n_136, wc5, n_117);
  not gc5 (wc5, n_120);
  or g122 (n_137, wc6, n_122);
  not gc6 (wc6, n_125);
  or g123 (n_45, wc7, n_99);
  not gc7 (wc7, n_100);
  or g124 (n_138, wc8, n_127);
  not gc8 (wc8, n_130);
  or g125 (n_106, wc9, n_102);
  not gc9 (wc9, n_103);
  or g126 (n_111, wc10, n_107);
  not gc10 (wc10, n_108);
  or g127 (n_116, wc11, n_112);
  not gc11 (wc11, n_113);
  or g128 (n_121, wc12, n_117);
  not gc12 (wc12, n_118);
  or g129 (n_126, wc13, n_122);
  not gc13 (wc13, n_123);
endmodule

module csa_tree_add_133_23_group_102_GENERIC(in_0, in_1, in_2, out_0);
  input [8:0] in_0, in_1, in_2;
  output [8:0] out_0;
  wire [8:0] in_0, in_1, in_2;
  wire [8:0] out_0;
  csa_tree_add_133_23_group_102_GENERIC_REAL g1(.in_0 (in_0), .in_1
       (in_1), .in_2 (in_2), .out_0 (out_0));
endmodule

module csa_tree_add_38_13_group_104_GENERIC_REAL(in_0, in_1, in_2,
     out_0);
// synthesis_equation "assign out_0 = ( $signed(in_2) + ( $signed(in_0) * $signed(in_1) )  )  ;"
  input [1:0] in_0;
  input [8:0] in_1;
  input [11:0] in_2;
  output [11:0] out_0;
  wire [1:0] in_0;
  wire [8:0] in_1;
  wire [11:0] in_2;
  wire [11:0] out_0;
  wire n_38, n_39, n_40, n_41, n_42, n_43, n_44, n_45;
  wire n_46, n_47, n_49, n_50, n_51, n_52, n_53, n_54;
  wire n_55, n_56, n_57, n_58, n_60, n_62, n_63, n_64;
  wire n_65, n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  wire n_73, n_74, n_76, n_77, n_79, n_85, n_86, n_87;
  wire n_88, n_89, n_90, n_91, n_92, n_93, n_94, n_95;
  wire n_96, n_97, n_98, n_99, n_100, n_101, n_102, n_103;
  wire n_104, n_105, n_106, n_107, n_108, n_109, n_110, n_111;
  wire n_112, n_113, n_114, n_115, n_116, n_117, n_121, n_123;
  wire n_126, n_127, n_128, n_129, n_131, n_132, n_133, n_134;
  wire n_136, n_137, n_138, n_140, n_141, n_142, n_143, n_145;
  wire n_146, n_147, n_148, n_150, n_151, n_152, n_153, n_155;
  wire n_156, n_157, n_158, n_160, n_161, n_162, n_163, n_165;
  wire n_166, n_167, n_168, n_170, n_171, n_172, n_173, n_175;
  wire n_176, n_177, n_178, n_179, n_180, n_181, n_182, n_183;
  wire n_184, n_185, n_186;
  and g2 (n_47, in_1[0], in_0[0]);
  and g3 (n_46, in_1[1], in_0[0]);
  and g4 (n_63, in_1[2], in_0[0]);
  and g5 (n_65, in_1[3], in_0[0]);
  and g6 (n_67, in_1[4], in_0[0]);
  and g7 (n_69, in_1[5], in_0[0]);
  and g8 (n_71, in_1[6], in_0[0]);
  and g9 (n_73, in_1[7], in_0[0]);
  nand g10 (n_76, in_1[8], in_0[0]);
  nand g11 (n_62, in_1[0], in_0[1]);
  nand g12 (n_64, in_1[1], in_0[1]);
  nand g13 (n_66, in_1[2], in_0[1]);
  nand g14 (n_68, in_1[3], in_0[1]);
  nand g15 (n_70, in_1[4], in_0[1]);
  nand g16 (n_72, in_1[5], in_0[1]);
  nand g17 (n_74, in_1[6], in_0[1]);
  nand g18 (n_77, in_1[7], in_0[1]);
  and g19 (n_79, in_1[8], in_0[1]);
  nand g35 (n_85, in_2[1], n_62);
  xor g37 (n_86, in_2[2], n_63);
  xor g38 (n_57, n_86, n_64);
  nand g39 (n_87, in_2[2], n_63);
  nand g40 (n_88, n_64, n_63);
  nand g41 (n_89, in_2[2], n_64);
  nand g42 (n_44, n_87, n_88, n_89);
  xor g43 (n_90, in_2[3], n_65);
  xor g44 (n_56, n_90, n_66);
  nand g45 (n_91, in_2[3], n_65);
  nand g46 (n_92, n_66, n_65);
  nand g47 (n_93, in_2[3], n_66);
  nand g48 (n_43, n_91, n_92, n_93);
  xor g49 (n_94, in_2[4], n_67);
  xor g50 (n_55, n_94, n_68);
  nand g51 (n_95, in_2[4], n_67);
  nand g52 (n_96, n_68, n_67);
  nand g53 (n_97, in_2[4], n_68);
  nand g54 (n_42, n_95, n_96, n_97);
  xor g55 (n_98, in_2[5], n_69);
  xor g56 (n_54, n_98, n_70);
  nand g57 (n_99, in_2[5], n_69);
  nand g58 (n_100, n_70, n_69);
  nand g59 (n_101, in_2[5], n_70);
  nand g60 (n_41, n_99, n_100, n_101);
  xor g61 (n_102, in_2[6], n_71);
  xor g62 (n_53, n_102, n_72);
  nand g63 (n_103, in_2[6], n_71);
  nand g64 (n_104, n_72, n_71);
  nand g65 (n_105, in_2[6], n_72);
  nand g66 (n_40, n_103, n_104, n_105);
  xor g67 (n_106, in_2[7], n_73);
  xor g68 (n_52, n_106, n_74);
  nand g69 (n_107, in_2[7], n_73);
  nand g70 (n_108, n_74, n_73);
  nand g71 (n_109, in_2[7], n_74);
  nand g72 (n_39, n_107, n_108, n_109);
  xor g75 (n_110, n_76, n_77);
  nand g77 (n_111, n_76, n_77);
  nand g80 (n_38, n_111, n_112, n_113);
  xor g81 (n_114, in_2[9], n_79);
  xor g82 (n_50, n_114, in_2[8]);
  nand g83 (n_115, in_2[9], n_79);
  nand g84 (n_116, in_2[8], n_79);
  nand g85 (n_117, in_2[9], in_2[8]);
  nand g86 (n_49, n_115, n_116, n_117);
  nand g93 (n_121, n_47, in_2[0]);
  nor g96 (n_123, n_46, n_58);
  nand g97 (n_126, n_46, n_58);
  nor g98 (n_128, n_45, n_57);
  nand g99 (n_131, n_45, n_57);
  nor g100 (n_133, n_44, n_56);
  nand g101 (n_136, n_44, n_56);
  nor g102 (n_60, n_43, n_55);
  nand g103 (n_140, n_43, n_55);
  nor g104 (n_142, n_42, n_54);
  nand g105 (n_145, n_42, n_54);
  nor g106 (n_147, n_41, n_53);
  nand g20 (n_150, n_41, n_53);
  nor g21 (n_152, n_40, n_52);
  nand g22 (n_155, n_40, n_52);
  nor g23 (n_157, n_39, n_51);
  nand g24 (n_160, n_39, n_51);
  nor g25 (n_162, n_38, n_50);
  nand g26 (n_165, n_38, n_50);
  nand g109 (n_129, n_126, n_127);
  nand g112 (n_134, n_131, n_132);
  nand g115 (n_138, n_136, n_137);
  nand g118 (n_143, n_140, n_141);
  nand g121 (n_148, n_145, n_146);
  nand g124 (n_153, n_150, n_151);
  nand g127 (n_158, n_155, n_156);
  nand g130 (n_163, n_160, n_161);
  nand g133 (n_168, n_165, n_166);
  nand g136 (n_173, n_170, n_171);
  xnor g141 (out_0[2], n_129, n_177);
  xnor g143 (out_0[3], n_134, n_178);
  xnor g145 (out_0[4], n_138, n_179);
  xnor g147 (out_0[5], n_143, n_180);
  xnor g149 (out_0[6], n_148, n_181);
  xnor g151 (out_0[7], n_153, n_182);
  xnor g153 (out_0[8], n_158, n_183);
  xnor g155 (out_0[9], n_163, n_184);
  xnor g157 (out_0[10], n_168, n_185);
  xnor g159 (out_0[11], n_173, n_186);
  xor g160 (out_0[0], in_2[0], n_47);
  xnor g164 (n_58, n_62, in_2[1]);
  or g166 (n_112, in_2[8], wc);
  not gc (wc, n_77);
  or g167 (n_113, in_2[8], wc0);
  not gc0 (wc0, n_76);
  or g168 (n_45, in_2[1], wc1, n_62);
  not gc1 (wc1, n_85);
  xnor g169 (n_51, n_110, in_2[8]);
  and g171 (n_172, in_2[10], wc2);
  not gc2 (wc2, in_2[11]);
  or g172 (n_175, in_2[10], wc3);
  not gc3 (wc3, in_2[11]);
  and g173 (n_167, in_2[10], wc4);
  not gc4 (wc4, n_49);
  or g174 (n_170, in_2[10], wc5);
  not gc5 (wc5, n_49);
  or g175 (n_127, n_121, n_123);
  or g176 (n_176, wc6, n_123);
  not gc6 (wc6, n_126);
  or g177 (n_186, wc7, n_172);
  not gc7 (wc7, n_175);
  xor g178 (out_0[1], n_121, n_176);
  or g179 (n_177, wc8, n_128);
  not gc8 (wc8, n_131);
  or g180 (n_178, wc9, n_133);
  not gc9 (wc9, n_136);
  or g181 (n_179, wc10, n_60);
  not gc10 (wc10, n_140);
  or g182 (n_180, wc11, n_142);
  not gc11 (wc11, n_145);
  or g183 (n_181, wc12, n_147);
  not gc12 (wc12, n_150);
  or g184 (n_182, wc13, n_152);
  not gc13 (wc13, n_155);
  or g185 (n_183, wc14, n_157);
  not gc14 (wc14, n_160);
  or g186 (n_184, wc15, n_162);
  not gc15 (wc15, n_165);
  or g187 (n_185, wc16, n_167);
  not gc16 (wc16, n_170);
  or g188 (n_132, wc17, n_128);
  not gc17 (wc17, n_129);
  or g189 (n_137, wc18, n_133);
  not gc18 (wc18, n_134);
  or g190 (n_141, wc19, n_60);
  not gc19 (wc19, n_138);
  or g191 (n_146, wc20, n_142);
  not gc20 (wc20, n_143);
  or g192 (n_151, wc21, n_147);
  not gc21 (wc21, n_148);
  or g193 (n_156, wc22, n_152);
  not gc22 (wc22, n_153);
  or g194 (n_161, wc23, n_157);
  not gc23 (wc23, n_158);
  or g195 (n_166, wc24, n_162);
  not gc24 (wc24, n_163);
  or g196 (n_171, n_167, wc25);
  not gc25 (wc25, n_168);
endmodule

module csa_tree_add_38_13_group_104_GENERIC(in_0, in_1, in_2, out_0);
  input [1:0] in_0;
  input [8:0] in_1;
  input [11:0] in_2;
  output [11:0] out_0;
  wire [1:0] in_0;
  wire [8:0] in_1;
  wire [11:0] in_2;
  wire [11:0] out_0;
  csa_tree_add_38_13_group_104_GENERIC_REAL g1(.in_0 (in_0), .in_1
       (in_1), .in_2 (in_2), .out_0 (out_0));
endmodule

module csa_tree_add_38_13_group_104_168_GENERIC_REAL(in_0, in_1, in_2,
     out_0);
// synthesis_equation "assign out_0 = ( $signed(in_2) + ( $signed(in_0) * $signed(in_1) )  )  ;"
  input [1:0] in_0;
  input [8:0] in_1;
  input [11:0] in_2;
  output [11:0] out_0;
  wire [1:0] in_0;
  wire [8:0] in_1;
  wire [11:0] in_2;
  wire [11:0] out_0;
  wire n_38, n_39, n_40, n_41, n_42, n_43, n_44, n_45;
  wire n_46, n_47, n_49, n_50, n_51, n_52, n_53, n_54;
  wire n_55, n_56, n_57, n_58, n_60, n_62, n_63, n_64;
  wire n_65, n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  wire n_73, n_74, n_76, n_77, n_79, n_85, n_86, n_87;
  wire n_88, n_89, n_90, n_91, n_92, n_93, n_94, n_95;
  wire n_96, n_97, n_98, n_99, n_100, n_101, n_102, n_103;
  wire n_104, n_105, n_106, n_107, n_108, n_109, n_110, n_111;
  wire n_112, n_113, n_114, n_115, n_116, n_117, n_121, n_123;
  wire n_126, n_127, n_128, n_129, n_131, n_132, n_133, n_134;
  wire n_136, n_137, n_138, n_140, n_141, n_142, n_143, n_145;
  wire n_146, n_147, n_148, n_150, n_151, n_152, n_153, n_155;
  wire n_156, n_157, n_158, n_160, n_161, n_162, n_163, n_165;
  wire n_166, n_167, n_168, n_170, n_171, n_172, n_173, n_175;
  wire n_176, n_177, n_178, n_179, n_180, n_181, n_182, n_183;
  wire n_184, n_185, n_186;
  and g2 (n_47, in_1[0], in_0[0]);
  and g3 (n_46, in_1[1], in_0[0]);
  and g4 (n_63, in_1[2], in_0[0]);
  and g5 (n_65, in_1[3], in_0[0]);
  and g6 (n_67, in_1[4], in_0[0]);
  and g7 (n_69, in_1[5], in_0[0]);
  and g8 (n_71, in_1[6], in_0[0]);
  and g9 (n_73, in_1[7], in_0[0]);
  nand g10 (n_76, in_1[8], in_0[0]);
  nand g11 (n_62, in_1[0], in_0[1]);
  nand g12 (n_64, in_1[1], in_0[1]);
  nand g13 (n_66, in_1[2], in_0[1]);
  nand g14 (n_68, in_1[3], in_0[1]);
  nand g15 (n_70, in_1[4], in_0[1]);
  nand g16 (n_72, in_1[5], in_0[1]);
  nand g17 (n_74, in_1[6], in_0[1]);
  nand g18 (n_77, in_1[7], in_0[1]);
  and g19 (n_79, in_1[8], in_0[1]);
  nand g35 (n_85, in_2[1], n_62);
  xor g37 (n_86, in_2[2], n_63);
  xor g38 (n_57, n_86, n_64);
  nand g39 (n_87, in_2[2], n_63);
  nand g40 (n_88, n_64, n_63);
  nand g41 (n_89, in_2[2], n_64);
  nand g42 (n_44, n_87, n_88, n_89);
  xor g43 (n_90, in_2[3], n_65);
  xor g44 (n_56, n_90, n_66);
  nand g45 (n_91, in_2[3], n_65);
  nand g46 (n_92, n_66, n_65);
  nand g47 (n_93, in_2[3], n_66);
  nand g48 (n_43, n_91, n_92, n_93);
  xor g49 (n_94, in_2[4], n_67);
  xor g50 (n_55, n_94, n_68);
  nand g51 (n_95, in_2[4], n_67);
  nand g52 (n_96, n_68, n_67);
  nand g53 (n_97, in_2[4], n_68);
  nand g54 (n_42, n_95, n_96, n_97);
  xor g55 (n_98, in_2[5], n_69);
  xor g56 (n_54, n_98, n_70);
  nand g57 (n_99, in_2[5], n_69);
  nand g58 (n_100, n_70, n_69);
  nand g59 (n_101, in_2[5], n_70);
  nand g60 (n_41, n_99, n_100, n_101);
  xor g61 (n_102, in_2[6], n_71);
  xor g62 (n_53, n_102, n_72);
  nand g63 (n_103, in_2[6], n_71);
  nand g64 (n_104, n_72, n_71);
  nand g65 (n_105, in_2[6], n_72);
  nand g66 (n_40, n_103, n_104, n_105);
  xor g67 (n_106, in_2[7], n_73);
  xor g68 (n_52, n_106, n_74);
  nand g69 (n_107, in_2[7], n_73);
  nand g70 (n_108, n_74, n_73);
  nand g71 (n_109, in_2[7], n_74);
  nand g72 (n_39, n_107, n_108, n_109);
  xor g75 (n_110, n_76, n_77);
  nand g77 (n_111, n_76, n_77);
  nand g80 (n_38, n_111, n_112, n_113);
  xor g81 (n_114, in_2[9], n_79);
  xor g82 (n_50, n_114, in_2[8]);
  nand g83 (n_115, in_2[9], n_79);
  nand g84 (n_116, in_2[8], n_79);
  nand g85 (n_117, in_2[9], in_2[8]);
  nand g86 (n_49, n_115, n_116, n_117);
  nand g93 (n_121, n_47, in_2[0]);
  nor g96 (n_123, n_46, n_58);
  nand g97 (n_126, n_46, n_58);
  nor g98 (n_128, n_45, n_57);
  nand g99 (n_131, n_45, n_57);
  nor g100 (n_133, n_44, n_56);
  nand g101 (n_136, n_44, n_56);
  nor g102 (n_60, n_43, n_55);
  nand g103 (n_140, n_43, n_55);
  nor g104 (n_142, n_42, n_54);
  nand g105 (n_145, n_42, n_54);
  nor g106 (n_147, n_41, n_53);
  nand g20 (n_150, n_41, n_53);
  nor g21 (n_152, n_40, n_52);
  nand g22 (n_155, n_40, n_52);
  nor g23 (n_157, n_39, n_51);
  nand g24 (n_160, n_39, n_51);
  nor g25 (n_162, n_38, n_50);
  nand g26 (n_165, n_38, n_50);
  nand g109 (n_129, n_126, n_127);
  nand g112 (n_134, n_131, n_132);
  nand g115 (n_138, n_136, n_137);
  nand g118 (n_143, n_140, n_141);
  nand g121 (n_148, n_145, n_146);
  nand g124 (n_153, n_150, n_151);
  nand g127 (n_158, n_155, n_156);
  nand g130 (n_163, n_160, n_161);
  nand g133 (n_168, n_165, n_166);
  nand g136 (n_173, n_170, n_171);
  xnor g141 (out_0[2], n_129, n_177);
  xnor g143 (out_0[3], n_134, n_178);
  xnor g145 (out_0[4], n_138, n_179);
  xnor g147 (out_0[5], n_143, n_180);
  xnor g149 (out_0[6], n_148, n_181);
  xnor g151 (out_0[7], n_153, n_182);
  xnor g153 (out_0[8], n_158, n_183);
  xnor g155 (out_0[9], n_163, n_184);
  xnor g157 (out_0[10], n_168, n_185);
  xnor g159 (out_0[11], n_173, n_186);
  xor g160 (out_0[0], in_2[0], n_47);
  xnor g164 (n_58, n_62, in_2[1]);
  or g166 (n_112, in_2[8], wc);
  not gc (wc, n_77);
  or g167 (n_113, in_2[8], wc0);
  not gc0 (wc0, n_76);
  or g168 (n_45, in_2[1], wc1, n_62);
  not gc1 (wc1, n_85);
  xnor g169 (n_51, n_110, in_2[8]);
  and g171 (n_172, in_2[10], wc2);
  not gc2 (wc2, in_2[11]);
  or g172 (n_175, in_2[10], wc3);
  not gc3 (wc3, in_2[11]);
  and g173 (n_167, in_2[10], wc4);
  not gc4 (wc4, n_49);
  or g174 (n_170, in_2[10], wc5);
  not gc5 (wc5, n_49);
  or g175 (n_127, n_121, n_123);
  or g176 (n_176, wc6, n_123);
  not gc6 (wc6, n_126);
  or g177 (n_186, wc7, n_172);
  not gc7 (wc7, n_175);
  xor g178 (out_0[1], n_121, n_176);
  or g179 (n_177, wc8, n_128);
  not gc8 (wc8, n_131);
  or g180 (n_178, wc9, n_133);
  not gc9 (wc9, n_136);
  or g181 (n_179, wc10, n_60);
  not gc10 (wc10, n_140);
  or g182 (n_180, wc11, n_142);
  not gc11 (wc11, n_145);
  or g183 (n_181, wc12, n_147);
  not gc12 (wc12, n_150);
  or g184 (n_182, wc13, n_152);
  not gc13 (wc13, n_155);
  or g185 (n_183, wc14, n_157);
  not gc14 (wc14, n_160);
  or g186 (n_184, wc15, n_162);
  not gc15 (wc15, n_165);
  or g187 (n_185, wc16, n_167);
  not gc16 (wc16, n_170);
  or g188 (n_132, wc17, n_128);
  not gc17 (wc17, n_129);
  or g189 (n_137, wc18, n_133);
  not gc18 (wc18, n_134);
  or g190 (n_141, wc19, n_60);
  not gc19 (wc19, n_138);
  or g191 (n_146, wc20, n_142);
  not gc20 (wc20, n_143);
  or g192 (n_151, wc21, n_147);
  not gc21 (wc21, n_148);
  or g193 (n_156, wc22, n_152);
  not gc22 (wc22, n_153);
  or g194 (n_161, wc23, n_157);
  not gc23 (wc23, n_158);
  or g195 (n_166, wc24, n_162);
  not gc24 (wc24, n_163);
  or g196 (n_171, n_167, wc25);
  not gc25 (wc25, n_168);
endmodule

module csa_tree_add_38_13_group_104_168_GENERIC(in_0, in_1, in_2,
     out_0);
  input [1:0] in_0;
  input [8:0] in_1;
  input [11:0] in_2;
  output [11:0] out_0;
  wire [1:0] in_0;
  wire [8:0] in_1;
  wire [11:0] in_2;
  wire [11:0] out_0;
  csa_tree_add_38_13_group_104_168_GENERIC_REAL g1(.in_0 (in_0), .in_1
       (in_1), .in_2 (in_2), .out_0 (out_0));
endmodule

module csa_tree_add_38_13_group_104_169_GENERIC_REAL(in_0, in_1, in_2,
     out_0);
// synthesis_equation "assign out_0 = ( $signed(in_2) + ( $signed(in_0) * $signed(in_1) )  )  ;"
  input [1:0] in_0;
  input [8:0] in_1;
  input [11:0] in_2;
  output [11:0] out_0;
  wire [1:0] in_0;
  wire [8:0] in_1;
  wire [11:0] in_2;
  wire [11:0] out_0;
  wire n_38, n_39, n_40, n_41, n_42, n_43, n_44, n_45;
  wire n_46, n_47, n_49, n_50, n_51, n_52, n_53, n_54;
  wire n_55, n_56, n_57, n_58, n_60, n_62, n_63, n_64;
  wire n_65, n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  wire n_73, n_74, n_76, n_77, n_79, n_85, n_86, n_87;
  wire n_88, n_89, n_90, n_91, n_92, n_93, n_94, n_95;
  wire n_96, n_97, n_98, n_99, n_100, n_101, n_102, n_103;
  wire n_104, n_105, n_106, n_107, n_108, n_109, n_110, n_111;
  wire n_112, n_113, n_114, n_115, n_116, n_117, n_121, n_123;
  wire n_126, n_127, n_128, n_129, n_131, n_132, n_133, n_134;
  wire n_136, n_137, n_138, n_140, n_141, n_142, n_143, n_145;
  wire n_146, n_147, n_148, n_150, n_151, n_152, n_153, n_155;
  wire n_156, n_157, n_158, n_160, n_161, n_162, n_163, n_165;
  wire n_166, n_167, n_168, n_170, n_171, n_172, n_173, n_175;
  wire n_176, n_177, n_178, n_179, n_180, n_181, n_182, n_183;
  wire n_184, n_185, n_186;
  and g2 (n_47, in_1[0], in_0[0]);
  and g3 (n_46, in_1[1], in_0[0]);
  and g4 (n_63, in_1[2], in_0[0]);
  and g5 (n_65, in_1[3], in_0[0]);
  and g6 (n_67, in_1[4], in_0[0]);
  and g7 (n_69, in_1[5], in_0[0]);
  and g8 (n_71, in_1[6], in_0[0]);
  and g9 (n_73, in_1[7], in_0[0]);
  nand g10 (n_76, in_1[8], in_0[0]);
  nand g11 (n_62, in_1[0], in_0[1]);
  nand g12 (n_64, in_1[1], in_0[1]);
  nand g13 (n_66, in_1[2], in_0[1]);
  nand g14 (n_68, in_1[3], in_0[1]);
  nand g15 (n_70, in_1[4], in_0[1]);
  nand g16 (n_72, in_1[5], in_0[1]);
  nand g17 (n_74, in_1[6], in_0[1]);
  nand g18 (n_77, in_1[7], in_0[1]);
  and g19 (n_79, in_1[8], in_0[1]);
  nand g35 (n_85, in_2[1], n_62);
  xor g37 (n_86, in_2[2], n_63);
  xor g38 (n_57, n_86, n_64);
  nand g39 (n_87, in_2[2], n_63);
  nand g40 (n_88, n_64, n_63);
  nand g41 (n_89, in_2[2], n_64);
  nand g42 (n_44, n_87, n_88, n_89);
  xor g43 (n_90, in_2[3], n_65);
  xor g44 (n_56, n_90, n_66);
  nand g45 (n_91, in_2[3], n_65);
  nand g46 (n_92, n_66, n_65);
  nand g47 (n_93, in_2[3], n_66);
  nand g48 (n_43, n_91, n_92, n_93);
  xor g49 (n_94, in_2[4], n_67);
  xor g50 (n_55, n_94, n_68);
  nand g51 (n_95, in_2[4], n_67);
  nand g52 (n_96, n_68, n_67);
  nand g53 (n_97, in_2[4], n_68);
  nand g54 (n_42, n_95, n_96, n_97);
  xor g55 (n_98, in_2[5], n_69);
  xor g56 (n_54, n_98, n_70);
  nand g57 (n_99, in_2[5], n_69);
  nand g58 (n_100, n_70, n_69);
  nand g59 (n_101, in_2[5], n_70);
  nand g60 (n_41, n_99, n_100, n_101);
  xor g61 (n_102, in_2[6], n_71);
  xor g62 (n_53, n_102, n_72);
  nand g63 (n_103, in_2[6], n_71);
  nand g64 (n_104, n_72, n_71);
  nand g65 (n_105, in_2[6], n_72);
  nand g66 (n_40, n_103, n_104, n_105);
  xor g67 (n_106, in_2[7], n_73);
  xor g68 (n_52, n_106, n_74);
  nand g69 (n_107, in_2[7], n_73);
  nand g70 (n_108, n_74, n_73);
  nand g71 (n_109, in_2[7], n_74);
  nand g72 (n_39, n_107, n_108, n_109);
  xor g75 (n_110, n_76, n_77);
  nand g77 (n_111, n_76, n_77);
  nand g80 (n_38, n_111, n_112, n_113);
  xor g81 (n_114, in_2[9], n_79);
  xor g82 (n_50, n_114, in_2[8]);
  nand g83 (n_115, in_2[9], n_79);
  nand g84 (n_116, in_2[8], n_79);
  nand g85 (n_117, in_2[9], in_2[8]);
  nand g86 (n_49, n_115, n_116, n_117);
  nand g93 (n_121, n_47, in_2[0]);
  nor g96 (n_123, n_46, n_58);
  nand g97 (n_126, n_46, n_58);
  nor g98 (n_128, n_45, n_57);
  nand g99 (n_131, n_45, n_57);
  nor g100 (n_133, n_44, n_56);
  nand g101 (n_136, n_44, n_56);
  nor g102 (n_60, n_43, n_55);
  nand g103 (n_140, n_43, n_55);
  nor g104 (n_142, n_42, n_54);
  nand g105 (n_145, n_42, n_54);
  nor g106 (n_147, n_41, n_53);
  nand g20 (n_150, n_41, n_53);
  nor g21 (n_152, n_40, n_52);
  nand g22 (n_155, n_40, n_52);
  nor g23 (n_157, n_39, n_51);
  nand g24 (n_160, n_39, n_51);
  nor g25 (n_162, n_38, n_50);
  nand g26 (n_165, n_38, n_50);
  nand g109 (n_129, n_126, n_127);
  nand g112 (n_134, n_131, n_132);
  nand g115 (n_138, n_136, n_137);
  nand g118 (n_143, n_140, n_141);
  nand g121 (n_148, n_145, n_146);
  nand g124 (n_153, n_150, n_151);
  nand g127 (n_158, n_155, n_156);
  nand g130 (n_163, n_160, n_161);
  nand g133 (n_168, n_165, n_166);
  nand g136 (n_173, n_170, n_171);
  xnor g141 (out_0[2], n_129, n_177);
  xnor g143 (out_0[3], n_134, n_178);
  xnor g145 (out_0[4], n_138, n_179);
  xnor g147 (out_0[5], n_143, n_180);
  xnor g149 (out_0[6], n_148, n_181);
  xnor g151 (out_0[7], n_153, n_182);
  xnor g153 (out_0[8], n_158, n_183);
  xnor g155 (out_0[9], n_163, n_184);
  xnor g157 (out_0[10], n_168, n_185);
  xnor g159 (out_0[11], n_173, n_186);
  xor g160 (out_0[0], in_2[0], n_47);
  xnor g164 (n_58, n_62, in_2[1]);
  or g166 (n_112, in_2[8], wc);
  not gc (wc, n_77);
  or g167 (n_113, in_2[8], wc0);
  not gc0 (wc0, n_76);
  or g168 (n_45, in_2[1], wc1, n_62);
  not gc1 (wc1, n_85);
  xnor g169 (n_51, n_110, in_2[8]);
  and g171 (n_172, in_2[10], wc2);
  not gc2 (wc2, in_2[11]);
  or g172 (n_175, in_2[10], wc3);
  not gc3 (wc3, in_2[11]);
  and g173 (n_167, in_2[10], wc4);
  not gc4 (wc4, n_49);
  or g174 (n_170, in_2[10], wc5);
  not gc5 (wc5, n_49);
  or g175 (n_127, n_121, n_123);
  or g176 (n_176, wc6, n_123);
  not gc6 (wc6, n_126);
  or g177 (n_186, wc7, n_172);
  not gc7 (wc7, n_175);
  xor g178 (out_0[1], n_121, n_176);
  or g179 (n_177, wc8, n_128);
  not gc8 (wc8, n_131);
  or g180 (n_178, wc9, n_133);
  not gc9 (wc9, n_136);
  or g181 (n_179, wc10, n_60);
  not gc10 (wc10, n_140);
  or g182 (n_180, wc11, n_142);
  not gc11 (wc11, n_145);
  or g183 (n_181, wc12, n_147);
  not gc12 (wc12, n_150);
  or g184 (n_182, wc13, n_152);
  not gc13 (wc13, n_155);
  or g185 (n_183, wc14, n_157);
  not gc14 (wc14, n_160);
  or g186 (n_184, wc15, n_162);
  not gc15 (wc15, n_165);
  or g187 (n_185, wc16, n_167);
  not gc16 (wc16, n_170);
  or g188 (n_132, wc17, n_128);
  not gc17 (wc17, n_129);
  or g189 (n_137, wc18, n_133);
  not gc18 (wc18, n_134);
  or g190 (n_141, wc19, n_60);
  not gc19 (wc19, n_138);
  or g191 (n_146, wc20, n_142);
  not gc20 (wc20, n_143);
  or g192 (n_151, wc21, n_147);
  not gc21 (wc21, n_148);
  or g193 (n_156, wc22, n_152);
  not gc22 (wc22, n_153);
  or g194 (n_161, wc23, n_157);
  not gc23 (wc23, n_158);
  or g195 (n_166, wc24, n_162);
  not gc24 (wc24, n_163);
  or g196 (n_171, n_167, wc25);
  not gc25 (wc25, n_168);
endmodule

module csa_tree_add_38_13_group_104_169_GENERIC(in_0, in_1, in_2,
     out_0);
  input [1:0] in_0;
  input [8:0] in_1;
  input [11:0] in_2;
  output [11:0] out_0;
  wire [1:0] in_0;
  wire [8:0] in_1;
  wire [11:0] in_2;
  wire [11:0] out_0;
  csa_tree_add_38_13_group_104_169_GENERIC_REAL g1(.in_0 (in_0), .in_1
       (in_1), .in_2 (in_2), .out_0 (out_0));
endmodule

